* NGSPICE file created from pll_3bitDiv.ext - technology: ihp-sg13g2

.subckt PLL_3BIT_DIV_PEX CLK_IN CLK_OUT Y0 Y2 Y1 VDD VSS nEN X1 X2 X0
X0 VDD a_53968_20434# a_53899_20488# VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0.19p ps=1.38u w=1u l=0.13u
X1 VSS 3bit_freq_divider_1.dff_nclk_0.nCLK a_61488_20220# VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=50.4f ps=0.66u w=0.42u l=0.13u
X2 a_62119_20605# a_61691_20534# a_61394_20220# VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0.1428p ps=1.52u w=0.42u l=0.13u
X3 a_52924_22885# 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.Q VDD VDD sg13_lv_pmos ad=0.3808p pd=2.92u as=0.2128p ps=1.5u w=1.12u l=0.13u
X4 a_53065_20179# a_53738_20514# a_53702_20612# VDD sg13_lv_pmos ad=0.17695p pd=1.56u as=43.05f ps=0.625u w=0.42u l=0.13u
X5 a_62119_22361# 3bit_freq_divider_1.dff_nclk_0.nCLK VDD VDD sg13_lv_pmos ad=0.1533p pd=1.57u as=0.11785p ps=1.025u w=0.42u l=0.13u
X6 a_53152_43159# VSS cap_cmim l=6.99u w=6.99u
X7 VDD a_52950_22157# 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.Q VDD sg13_lv_pmos ad=0.2016p pd=1.5u as=0.3808p ps=2.92u w=1.12u l=0.13u
X8 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 3bit_freq_divider_1.sg13g2_nand2_1_0.Y VSS VSS sg13_lv_nmos ad=0.259p pd=2.18u as=0.259p ps=2.18u w=0.74u l=0.13u
X9 VSS 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.Q a_61061_23234# VSS sg13_lv_nmos ad=0.1331p pd=1.12u as=0.1216p ps=1.02u w=0.64u l=0.13u
X10 a_62879_24125# a_61887_24046# a_62654_23727# VDD sg13_lv_pmos ad=43.05f pd=0.625u as=0.17695p ps=1.56u w=0.42u l=0.13u
X11 a_53022_43738# a_53022_43738# VDD VDD sg13_lv_pmos ad=59f pd=0.74u as=0.104p ps=1.34u w=0.2u l=0.13u
X12 VSS a_55345_24897# 3bit_freq_divider_0.freq_div_cell_0.Cin VSS sg13_lv_nmos ad=0.1331p pd=1.12u as=0.2516p ps=2.16u w=0.74u l=0.13u
X13 a_64383_23434# a_64383_23628# VSS VSS sg13_lv_nmos ad=0.2516p pd=2.16u as=0.1544p ps=1.235u w=0.74u l=0.13u
X14 VDD a_53774_21934# a_53738_22270# VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0.34p ps=2.68u w=1u l=0.13u
X15 a_55485_23233# 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.Q VSS VSS sg13_lv_nmos ad=0.1216p pd=1.02u as=0.1331p ps=1.12u w=0.64u l=0.13u
X16 a_64383_23300# a_64383_23628# a_64424_22200# VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0.1428p ps=1.52u w=0.42u l=0.13u
X17 VSS charge_pump_0.vout VSS VSS sg13_lv_nmos ad=0.285p pd=1.88u as=0.53383n ps=1.58949m w=1.5u l=0.65u
X18 VDD a_53022_43738# a_57084_43159# VDD sg13_lv_pmos ad=0.104p pd=1.34u as=59f ps=0.74u w=0.2u l=0.13u
X19 VDD a_51648_21103# 3bit_freq_divider_0.dff_nclk_0.nCLK VDD sg13_lv_pmos ad=0.3822p pd=1.84u as=0.3808p ps=2.92u w=1.12u l=0.13u
X20 a_64383_23434# a_64383_23628# VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0.19p ps=1.38u w=1u l=0.13u
X21 a_54627_42591# vco_wob_0.vctl VSS VSS sg13_lv_nmos ad=65.99999f pd=0.74u as=0.102p ps=1.28u w=0.3u l=0.13u
X22 a_59799_40285# 3bit_freq_divider_0.CLK_IN a_58515_40413# VDD sg13_lv_pmos ad=0.17p pd=1.68u as=0.1106p ps=0.945u w=0.5u l=0.13u
X23 a_61972_23244# 3bit_freq_divider_1.freq_div_cell_0.Cin VSS VSS sg13_lv_nmos ad=88.8f pd=0.98u as=0.15245p ps=1.17u w=0.74u l=0.13u
X24 a_54494_43159# a_53152_43159# a_54627_42591# VSS sg13_lv_nmos ad=0.11p pd=0.94u as=0.17p ps=1.68u w=0.5u l=0.13u
X25 a_54427_40283# a_54489_40413# a_53147_40413# VDD sg13_lv_pmos ad=0.11p pd=0.94u as=0.11p ps=0.94u w=0.5u l=0.13u
X26 VDD 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.D a_54504_23771# VDD sg13_lv_pmos ad=0.1428p pd=1.52u as=79.8f ps=0.8u w=0.42u l=0.13u
X27 a_53774_20178# 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.sg13g2_dfrbp_1_0.CLK VSS VSS sg13_lv_nmos ad=0.2516p pd=2.16u as=0.1544p ps=1.235u w=0.74u l=0.13u
X28 a_54504_20259# 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.D a_55086_20219# VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=50.4f ps=0.66u w=0.42u l=0.13u
X29 charge_pump_0.bias_n charge_pump_0.bias_n VSS VSS sg13_lv_nmos ad=0.34p pd=2.68u as=0.34p ps=2.68u w=1u l=1u
X30 VSS 3bit_freq_divider_0.freq_div_cell_0.Cout a_54434_21392# VSS sg13_lv_nmos ad=0.374p pd=2.46u as=0.17462p ps=1.185u w=0.55u l=0.13u
X31 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.Q a_63463_23728# VSS VSS sg13_lv_nmos ad=0.2516p pd=2.16u as=0.14505p ps=1.15u w=0.74u l=0.13u
X32 a_47954_28913# PFD_0.VCO_CLK a_48909_28913# VSS sg13_lv_nmos ad=68.39999f pd=0.74u as=68.39999f ps=0.74u w=0.36u l=0.15u
X33 a_54898_21129# 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.Q a_54434_21392# VDD sg13_lv_pmos ad=0.1225p pd=1.245u as=0.34p ps=2.68u w=1u l=0.13u
X34 VSS charge_pump_0.vout VSS VSS sg13_lv_nmos ad=0.285p pd=1.88u as=0 ps=0 w=1.5u l=0.65u
X35 a_51693_23426# 3bit_freq_divider_0.dff_nclk_0.nRST VDD VDD sg13_lv_pmos ad=0.1533p pd=1.57u as=0.11785p ps=1.025u w=0.42u l=0.13u
X36 3bit_freq_divider_1.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 3bit_freq_divider_1.dff_nclk_0.nCLK VSS VSS sg13_lv_nmos ad=0.259p pd=2.18u as=0.259p ps=2.18u w=0.74u l=0.13u
X37 PFD_0.UP a_47777_29803# VSS VSS sg13_lv_nmos ad=0.1632p pd=1.64u as=0.1632p ps=1.64u w=0.48u l=0.15u
X38 VDD a_62654_23727# a_62900_23691# VDD sg13_lv_pmos ad=0.2163p pd=1.55u as=79.8f ps=0.8u w=0.42u l=0.13u
X39 a_54504_23771# 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.D a_55086_23731# VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=50.4f ps=0.66u w=0.42u l=0.13u
X40 a_60967_23234# 3bit_freq_divider_1.freq_div_cell_0.Cin VDD VDD sg13_lv_pmos ad=0.1596p pd=1.22u as=0.2856p ps=2.36u w=0.84u l=0.13u
X41 a_54602_23243# 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.Q 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.D VSS sg13_lv_nmos ad=88.8f pd=0.98u as=0.1628p ps=1.18u w=0.74u l=0.13u
X42 a_54898_24641# 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.Q a_54434_24904# VDD sg13_lv_pmos ad=0.1225p pd=1.245u as=0.34p ps=2.68u w=1u l=0.13u
X43 VDD 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.Q a_60967_21478# VDD sg13_lv_pmos ad=0.1918p pd=1.5u as=0.1596p ps=1.22u w=0.84u l=0.13u
X44 a_62221_24117# a_61691_24046# a_62119_24117# VDD sg13_lv_pmos ad=51.45f pd=0.665u as=79.8f ps=0.8u w=0.42u l=0.13u
X45 a_58426_43159# a_57178_43159# 3bit_freq_divider_0.CLK_IN VDD sg13_lv_pmos ad=0.11p pd=0.94u as=0.1106p ps=0.945u w=0.5u l=0.13u
X46 a_62246_20260# a_61887_20534# a_62119_20605# VSS sg13_lv_nmos ad=54.6f pd=0.68u as=79.8f ps=0.8u w=0.42u l=0.13u
X47 a_52074_23051# a_51684_22692# a_51693_23426# VSS sg13_lv_nmos ad=54.6f pd=0.68u as=79.8f ps=0.8u w=0.42u l=0.13u
X48 a_54504_22015# 3bit_freq_divider_0.dff_nclk_0.nCLK VDD VDD sg13_lv_pmos ad=79.8f pd=0.8u as=0.1428p ps=1.52u w=0.42u l=0.13u
X49 VDD a_55345_23141# 3bit_freq_divider_0.freq_div_cell_0.Cout VDD sg13_lv_pmos ad=0.1918p pd=1.5u as=0.3808p ps=2.92u w=1.12u l=0.13u
X50 a_64464_23130# a_64419_23326# a_64464_23052# VSS sg13_lv_nmos ad=48.3f pd=0.65u as=54.6f ps=0.68u w=0.42u l=0.13u
X51 VSS a_63255_21488# 3bit_freq_divider_1.sg13g2_or3_1_0.A VSS sg13_lv_nmos ad=0.3108p pd=2.32u as=0.1628p ps=1.18u w=0.74u l=0.13u
X52 a_61675_22886# 3bit_freq_divider_1.freq_div_cell_0.Cin VDD VDD sg13_lv_pmos ad=0.1225p pd=1.245u as=0.36p ps=2.72u w=1u l=0.13u
X53 VDD a_53022_43738# a_53085_40283# VDD sg13_lv_pmos ad=0.104p pd=1.34u as=59.75f ps=0.745u w=0.2u l=0.13u
X54 a_53968_20434# a_53738_20514# a_54324_20259# VSS sg13_lv_nmos ad=79.8f pd=0.8u as=54.6f ps=0.68u w=0.42u l=0.13u
X55 VSS 3bit_freq_divider_0.sg13g2_or3_1_0.B a_51648_21103# VSS sg13_lv_nmos ad=0.1045p pd=0.93u as=0.198p ps=1.27u w=0.55u l=0.13u
X56 VDD 3bit_freq_divider_0.EN charge_pump_0.bias_p VDD sg13_lv_pmos ad=0.17p pd=1.68u as=0.17p ps=1.68u w=0.5u l=0.15u
X57 a_55345_23141# 3bit_freq_divider_0.freq_div_cell_0.Cin a_55485_23233# VSS sg13_lv_nmos ad=0.2176p pd=1.96u as=0.1216p ps=1.02u w=0.64u l=0.13u
X58 charge_pump_0.bias_n charge_pump_0.bias_p a_55862_56737# VDD sg13_lv_pmos ad=0.68p pd=4.68u as=0.38p ps=2.38u w=2u l=1u
X59 a_53152_43159# a_52944_43077# a_53058_43159# VDD sg13_lv_pmos ad=0.1106p pd=0.945u as=0.17p ps=1.68u w=0.5u l=0.13u
X60 VDD a_53022_43738# a_55769_40283# VDD sg13_lv_pmos ad=59f pd=0.74u as=59f ps=0.74u w=0.2u l=0.13u
X61 3bit_freq_divider_1.sg13g2_tiehi_1.L_HI a_60584_24580# a_60385_24558# VDD sg13_lv_pmos ad=0.3927p pd=2.99u as=0.4657p ps=2.54u w=1.155u l=0.13u
X62 a_54324_20259# a_53899_20488# a_54252_20259# VSS sg13_lv_nmos ad=54.6f pd=0.68u as=48.3f ps=0.65u w=0.42u l=0.13u
X63 a_62270_24055# a_62119_24117# VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0.34p ps=2.68u w=1u l=0.13u
X64 a_62324_22016# a_62270_22299# a_62246_22016# VSS sg13_lv_nmos ad=48.3f pd=0.65u as=54.6f ps=0.68u w=0.42u l=0.13u
X65 VDD X2 a_52924_21129# VDD sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X66 a_52944_43077# a_53147_40413# a_53085_40283# VDD sg13_lv_pmos ad=0.11p pd=0.94u as=0.17p ps=1.68u w=0.5u l=0.13u
X67 VSS a_53774_21934# a_53738_22270# VSS sg13_lv_nmos ad=0.1544p pd=1.235u as=0.2516p ps=2.16u w=0.74u l=0.13u
X68 a_46749_30782# CLK_IN a_45579_29803# VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=79.8f ps=0.8u w=0.42u l=0.15u
X69 a_54400_43159# a_53152_43159# a_54494_43159# VDD sg13_lv_pmos ad=0.11p pd=0.94u as=0.1106p ps=0.945u w=0.5u l=0.13u
X70 3bit_freq_divider_1.freq_div_cell_0.Cin a_60967_24990# VDD VDD sg13_lv_pmos ad=0.3808p pd=2.92u as=0.1918p ps=1.5u w=1.12u l=0.13u
X71 a_55742_43159# a_53022_43738# VDD VDD sg13_lv_pmos ad=59.75f pd=0.745u as=0.104p ps=1.34u w=0.2u l=0.13u
X72 a_53968_23946# a_53738_24026# a_54324_23771# VSS sg13_lv_nmos ad=79.8f pd=0.8u as=54.6f ps=0.68u w=0.42u l=0.13u
X73 a_63038_20215# 3bit_freq_divider_1.dff_nclk_0.nCLK VSS VSS sg13_lv_nmos ad=47.25f pd=0.645u as=90.3f ps=0.85u w=0.42u l=0.13u
X74 a_62900_20179# a_62654_20215# a_63038_20215# VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=47.25f ps=0.645u w=0.42u l=0.13u
X75 3bit_freq_divider_0.sg13g2_or3_1_0.C a_52886_24904# VSS VSS sg13_lv_nmos ad=0.1628p pd=1.18u as=0.3108p ps=2.32u w=0.74u l=0.13u
X76 VDD a_53022_43738# a_57111_40283# VDD sg13_lv_pmos ad=59f pd=0.74u as=59f ps=0.74u w=0.2u l=0.13u
X77 a_48909_28913# PFD_0.VCO_CLK a_47954_28913# VSS sg13_lv_nmos ad=0.1224p pd=1.4u as=68.39999f ps=0.74u w=0.36u l=0.15u
X78 a_54324_23771# a_53899_24000# a_54252_23771# VSS sg13_lv_nmos ad=54.6f pd=0.68u as=48.3f ps=0.65u w=0.42u l=0.13u
X79 VSS vco_wob_0.vctl a_58454_40850# VSS sg13_lv_nmos ad=0.102p pd=1.28u as=65.99999f ps=0.74u w=0.3u l=0.13u
X80 a_58453_40283# a_53022_43738# VDD VDD sg13_lv_pmos ad=59f pd=0.74u as=0.104p ps=1.34u w=0.2u l=0.13u
X81 a_53899_22244# a_53774_21934# a_53065_21935# VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0.17695p ps=1.56u w=1u l=0.13u
X82 VDD X0 a_52924_24641# VDD sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X83 VDD a_64384_21091# 3bit_freq_divider_1.dff_nclk_0.nCLK VDD sg13_lv_pmos ad=0.3822p pd=1.84u as=0.3808p ps=2.92u w=1.12u l=0.13u
X84 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.D 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.Q a_61972_23244# VSS sg13_lv_nmos ad=0.1628p pd=1.18u as=88.8f ps=0.98u w=0.74u l=0.13u
X85 VDD 3bit_freq_divider_1.sg13g2_tiehi_1.L_HI a_61878_24642# VDD sg13_lv_pmos ad=0.2128p pd=1.5u as=0.3808p ps=2.92u w=1.12u l=0.13u
X86 3bit_freq_divider_1.sg13g2_or3_1_0.B a_63255_23244# a_63426_22886# VDD sg13_lv_pmos ad=0.3808p pd=2.92u as=0.2128p ps=1.5u w=1.12u l=0.13u
X87 VSS vco_wob_0.vctl a_53022_43738# VSS sg13_lv_nmos ad=0.102p pd=1.28u as=65.99999f ps=0.74u w=0.3u l=0.13u
X88 a_51729_23026# a_51631_22774# a_51693_23426# VDD sg13_lv_pmos ad=51.45f pd=0.665u as=79.8f ps=0.8u w=0.42u l=0.13u
X89 a_53147_40413# VSS cap_cmim l=6.99u w=6.99u
X90 a_57084_43159# a_53022_43738# VDD VDD sg13_lv_pmos ad=59.75f pd=0.745u as=0.104p ps=1.34u w=0.2u l=0.13u
X91 a_61887_20534# a_61691_20534# VSS VSS sg13_lv_nmos ad=0.2516p pd=2.16u as=0.1544p ps=1.235u w=0.74u l=0.13u
X92 a_54400_43159# a_53152_43159# a_54494_43159# VDD sg13_lv_pmos ad=0.17p pd=1.68u as=0.11p ps=0.94u w=0.5u l=0.13u
X93 a_62119_22361# a_61691_22290# a_61394_21976# VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0.1428p ps=1.52u w=0.42u l=0.13u
X94 a_52950_23913# a_53065_23691# VDD VDD sg13_lv_pmos ad=0.2856p pd=2.36u as=0.2016p ps=1.5u w=0.84u l=0.13u
X95 a_54504_20259# a_53738_20514# a_53968_20434# VDD sg13_lv_pmos ad=0.1428p pd=1.52u as=79.8f ps=0.8u w=0.42u l=0.13u
X96 a_62119_24117# 3bit_freq_divider_1.dff_nclk_0.nCLK VDD VDD sg13_lv_pmos ad=0.1533p pd=1.57u as=0.11785p ps=1.025u w=0.42u l=0.13u
X97 PFD_0.VCO_CLK PFD_0.VCO_CLK a_46817_27899# VDD sg13_lv_pmos ad=60.8f pd=0.7u as=0.1088p ps=1.32u w=0.32u l=0.15u
X98 VDD 3bit_freq_divider_0.CLK_IN 3bit_freq_divider_1.sg13g2_nand2_1_0.Y VDD sg13_lv_pmos ad=0.3808p pd=2.92u as=0.2128p ps=1.5u w=1.12u l=0.13u
X99 VDD a_62900_21935# a_62879_22369# VDD sg13_lv_pmos ad=79.8f pd=0.8u as=43.05f ps=0.625u w=0.42u l=0.13u
X100 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 3bit_freq_divider_1.sg13g2_nand2_1_0.Y VDD VDD sg13_lv_pmos ad=0.392p pd=2.94u as=0.392p ps=2.94u w=1.12u l=0.13u
X101 a_53350_21129# X2 a_52886_21392# VDD sg13_lv_pmos ad=0.1225p pd=1.245u as=0.34p ps=2.68u w=1u l=0.13u
X102 a_58454_40850# a_58515_40413# a_57173_40413# VSS sg13_lv_nmos ad=0.17p pd=1.68u as=0.11p ps=0.94u w=0.5u l=0.13u
X103 VSS 3bit_freq_divider_0.EN a_56055_21027# VSS sg13_lv_nmos ad=0.2516p pd=2.16u as=66.6f ps=0.92u w=0.74u l=0.13u
X104 VDD a_62654_23727# a_63463_23728# VDD sg13_lv_pmos ad=0.2016p pd=1.5u as=0.2856p ps=2.36u w=0.84u l=0.13u
X105 VSS charge_pump_0.vout VSS VSS sg13_lv_nmos ad=0.285p pd=1.88u as=0 ps=0 w=1.5u l=0.65u
X106 a_55742_43159# a_54494_43159# a_55836_43159# VDD sg13_lv_pmos ad=0.17p pd=1.68u as=0.11p ps=0.94u w=0.5u l=0.13u
X107 a_62654_21971# a_61887_22290# a_62270_22299# VSS sg13_lv_nmos ad=0.2017p pd=1.48u as=0.19397p ps=1.29u w=0.64u l=0.13u
X108 VSS a_62900_20179# a_62848_20215# VSS sg13_lv_nmos ad=90.3f pd=0.85u as=54.6f ps=0.68u w=0.42u l=0.13u
X109 VSS 3bit_freq_divider_0.sg13g2_nand2_1_0.Y 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK VSS sg13_lv_nmos ad=0.259p pd=2.18u as=0.259p ps=2.18u w=0.74u l=0.13u
X110 a_61394_23732# 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.D VDD VDD sg13_lv_pmos ad=79.8f pd=0.8u as=0.1428p ps=1.52u w=0.42u l=0.13u
X111 a_62848_20215# a_61691_20534# a_62654_20215# VSS sg13_lv_nmos ad=54.6f pd=0.68u as=0.2017p ps=1.48u w=0.42u l=0.13u
X112 a_53774_21934# 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK VSS VSS sg13_lv_nmos ad=0.2516p pd=2.16u as=0.1544p ps=1.235u w=0.74u l=0.13u
X113 a_53054_23243# X1 3bit_freq_divider_0.sg13g2_or3_1_0.B VSS sg13_lv_nmos ad=88.8f pd=0.98u as=0.1628p ps=1.18u w=0.74u l=0.13u
X114 a_53350_24641# X0 a_52886_24904# VDD sg13_lv_pmos ad=0.1225p pd=1.245u as=0.34p ps=2.68u w=1u l=0.13u
X115 VDD a_53022_43738# a_58426_43159# VDD sg13_lv_pmos ad=0.104p pd=1.34u as=59f ps=0.74u w=0.2u l=0.13u
X116 a_56038_24617# a_55941_24882# 3bit_freq_divider_0.sg13g2_tiehi_1.L_HI VDD sg13_lv_pmos ad=0.4657p pd=2.54u as=0.3927p ps=2.99u w=1.155u l=0.13u
X117 VDD 3bit_freq_divider_0.dff_nclk_0.nCLK a_53445_20214# VDD sg13_lv_pmos ad=79.8f pd=0.8u as=79.8f ps=0.8u w=0.42u l=0.13u
X118 VSS charge_pump_0.vout VSS VSS sg13_lv_nmos ad=0.285p pd=1.88u as=0 ps=0 w=1.5u l=0.65u
X119 a_57112_40850# vco_wob_0.vctl VSS VSS sg13_lv_nmos ad=65.99999f pd=0.74u as=0.102p ps=1.28u w=0.3u l=0.13u
X120 a_60584_24580# a_60385_24717# a_60479_25023# VSS sg13_lv_nmos ad=0.27427p pd=2.28u as=0.2307p ps=1.615u w=0.795u l=0.13u
X121 VSS a_61707_21488# 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.D VSS sg13_lv_nmos ad=0.3108p pd=2.32u as=0.1628p ps=1.18u w=0.74u l=0.13u
X122 a_63255_25000# Y0 a_63223_24642# VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0.1225p ps=1.245u w=1u l=0.13u
X123 VDD a_51648_24041# a_51685_23725# VDD sg13_lv_pmos ad=0.2163p pd=1.55u as=79.8f ps=0.8u w=0.42u l=0.13u
X124 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.Q a_63463_20216# VDD VDD sg13_lv_pmos ad=0.3808p pd=2.92u as=0.2016p ps=1.5u w=1.12u l=0.13u
X125 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.D a_54434_21392# VSS VSS sg13_lv_nmos ad=0.1628p pd=1.18u as=0.3108p ps=2.32u w=0.74u l=0.13u
X126 VSS Y0 a_63255_25000# VSS sg13_lv_nmos ad=0.15245p pd=1.17u as=0.17462p ps=1.185u w=0.55u l=0.13u
X127 VSS a_56887_49467# VSS VSS sg13_lv_nmos ad=95f pd=0.88u as=0 ps=0 w=0.5u l=0.65u
X128 a_48909_28913# PFD_0.VCO_CLK a_47954_28913# VSS sg13_lv_nmos ad=68.39999f pd=0.74u as=0.1224p ps=1.4u w=0.36u l=0.15u
X129 VDD a_62270_20543# a_62221_20605# VDD sg13_lv_pmos ad=0.11785p pd=1.025u as=51.45f ps=0.665u w=0.42u l=0.13u
X130 a_62246_22016# a_61887_22290# a_62119_22361# VSS sg13_lv_nmos ad=54.6f pd=0.68u as=79.8f ps=0.8u w=0.42u l=0.13u
X131 VDD 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.Q a_63426_21130# VDD sg13_lv_pmos ad=0.2128p pd=1.5u as=0.3808p ps=2.92u w=1.12u l=0.13u
X132 VDD 3bit_freq_divider_0.freq_div_cell_0.Cout a_54898_21129# VDD sg13_lv_pmos ad=0.36p pd=2.72u as=0.1225p ps=1.245u w=1u l=0.13u
X133 VSS charge_pump_0.vout VSS VSS sg13_lv_nmos ad=0.285p pd=1.88u as=0 ps=0 w=1.5u l=0.65u
X134 a_64362_24865# a_64459_24995# a_64731_24890# VDD sg13_lv_pmos ad=0.2442p pd=2.06u as=0.4657p ps=2.54u w=0.66u l=0.13u
X135 a_55831_40413# a_57173_40413# a_57112_40850# VSS sg13_lv_nmos ad=0.11p pd=0.94u as=0.17p ps=1.68u w=0.5u l=0.13u
X136 VSS a_56887_49467# VSS VSS sg13_lv_nmos ad=95f pd=0.88u as=0 ps=0 w=0.5u l=0.65u
X137 a_47777_29803# a_46749_30782# VSS VSS sg13_lv_nmos ad=0.1224p pd=1.4u as=0.1224p ps=1.4u w=0.36u l=0.15u
X138 a_55086_21975# 3bit_freq_divider_0.dff_nclk_0.nCLK VSS VSS sg13_lv_nmos ad=50.4f pd=0.66u as=0.1428p ps=1.52u w=0.42u l=0.13u
X139 VDD 3bit_freq_divider_0.sg13g2_tiehi_1.L_HI a_54898_24641# VDD sg13_lv_pmos ad=0.36p pd=2.72u as=0.1225p ps=1.245u w=1u l=0.13u
X140 a_53445_21970# a_53065_21935# VDD VDD sg13_lv_pmos ad=79.8f pd=0.8u as=0.2163p ps=1.55u w=0.42u l=0.13u
X141 VSS 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.Q a_52886_23148# VSS sg13_lv_nmos ad=0.374p pd=2.46u as=0.17462p ps=1.185u w=0.55u l=0.13u
X142 a_64384_21091# 3bit_freq_divider_1.sg13g2_or3_1_0.A VSS VSS sg13_lv_nmos ad=0.198p pd=1.27u as=0.13395p ps=1.12u w=0.55u l=0.13u
X143 a_63255_23244# 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.Q VSS VSS sg13_lv_nmos ad=0.17462p pd=1.185u as=0.374p ps=2.46u w=0.55u l=0.13u
X144 a_54494_43159# a_53152_43159# a_54400_43159# VDD sg13_lv_pmos ad=0.1106p pd=0.945u as=0.17p ps=1.68u w=0.5u l=0.13u
X145 a_63426_24642# Y0 VDD VDD sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X146 a_62270_20543# a_62119_20605# VSS VSS sg13_lv_nmos ad=0.19397p pd=1.29u as=0.1825p ps=1.325u w=0.64u l=0.13u
X147 VSS a_56887_49467# VSS VSS sg13_lv_nmos ad=95f pd=0.88u as=0 ps=0 w=0.5u l=0.65u
X148 VSS vco_wob_0.vctl a_58653_42591# VSS sg13_lv_nmos ad=0.102p pd=1.28u as=65.99999f ps=0.74u w=0.3u l=0.13u
X149 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.nQ a_62654_21971# VSS VSS sg13_lv_nmos ad=0.2775p pd=2.23u as=0.2516p ps=2.16u w=0.74u l=0.13u
X150 a_58653_42591# a_57178_43159# 3bit_freq_divider_0.CLK_IN VSS sg13_lv_nmos ad=0.17p pd=1.68u as=0.11p ps=0.94u w=0.5u l=0.13u
X151 VDD a_64383_23889# a_64384_24445# VDD sg13_lv_pmos ad=0.2016p pd=1.5u as=0.2856p ps=2.36u w=0.84u l=0.13u
X152 a_51708_21299# 3bit_freq_divider_0.sg13g2_or3_1_0.A VDD VDD sg13_lv_pmos ad=0.22p pd=1.44u as=0.3822p ps=1.84u w=1u l=0.13u
X153 VSS 3bit_freq_divider_0.dff_nclk_0.nRST a_52074_23129# VSS sg13_lv_nmos ad=0.1825p pd=1.325u as=48.3f ps=0.65u w=0.42u l=0.13u
X154 a_53147_40413# a_54489_40413# a_54427_40283# VDD sg13_lv_pmos ad=0.11p pd=0.94u as=0.17p ps=1.68u w=0.5u l=0.13u
X155 VDD 3bit_freq_divider_0.sg13g2_nand2_1_0.Y 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.sg13g2_dfrbp_1_0.CLK VDD sg13_lv_pmos ad=0.392p pd=2.94u as=0.392p ps=2.94u w=1.12u l=0.13u
X156 a_57178_43159# VSS cap_cmim l=6.99u w=6.99u
X157 VSS charge_pump_0.vout VSS VSS sg13_lv_nmos ad=0.51p pd=3.68u as=0 ps=0 w=1.5u l=0.65u
X158 VSS charge_pump_0.vout VSS VSS sg13_lv_nmos ad=0.285p pd=1.88u as=0 ps=0 w=1.5u l=0.65u
X159 VSS a_56887_49467# VSS VSS sg13_lv_nmos ad=95f pd=0.88u as=0 ps=0 w=0.5u l=0.65u
X160 a_62879_20613# a_61887_20534# a_62654_20215# VDD sg13_lv_pmos ad=43.05f pd=0.625u as=0.17695p ps=1.56u w=0.42u l=0.13u
X161 a_61887_22290# a_61691_22290# VSS VSS sg13_lv_nmos ad=0.2516p pd=2.16u as=0.1544p ps=1.235u w=0.74u l=0.13u
X162 VSS a_52950_22157# 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.Q VSS sg13_lv_nmos ad=0.14505p pd=1.15u as=0.2516p ps=2.16u w=0.74u l=0.13u
X163 VSS a_56887_49467# VSS VSS sg13_lv_nmos ad=95f pd=0.88u as=0 ps=0 w=0.5u l=0.65u
X164 a_63520_25000# 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.Q VSS VSS sg13_lv_nmos ad=88.8f pd=0.98u as=0.15245p ps=1.17u w=0.74u l=0.13u
X165 a_53702_24124# a_53445_23726# VDD VDD sg13_lv_pmos ad=43.05f pd=0.625u as=79.8f ps=0.8u w=0.42u l=0.13u
X166 a_61707_25000# 3bit_freq_divider_1.sg13g2_tiehi_1.L_HI VSS VSS sg13_lv_nmos ad=0.17462p pd=1.185u as=0.374p ps=2.46u w=0.55u l=0.13u
X167 VDD 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK a_61691_22290# VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0.34p ps=2.68u w=1u l=0.13u
X168 VDD 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.Q a_54472_21129# VDD sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X169 VSS 3bit_freq_divider_0.freq_div_cell_0.Cin a_54602_23243# VSS sg13_lv_nmos ad=0.15245p pd=1.17u as=88.8f ps=0.98u w=0.74u l=0.13u
X170 VSS a_51648_24041# a_51648_24438# VSS sg13_lv_nmos ad=0.14505p pd=1.15u as=0.187p ps=1.78u w=0.55u l=0.13u
X171 VSS charge_pump_0.vout VSS VSS sg13_lv_nmos ad=0.285p pd=1.88u as=0 ps=0 w=1.5u l=0.65u
X172 a_53147_40413# a_54489_40413# a_54427_40283# VDD sg13_lv_pmos ad=0.1106p pd=0.945u as=0.11p ps=0.94u w=0.5u l=0.13u
X173 a_62270_20543# a_62119_20605# VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0.34p ps=2.68u w=1u l=0.13u
X174 a_51648_21103# 3bit_freq_divider_0.sg13g2_or3_1_0.C a_51708_21413# VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0.1275p ps=1.255u w=1u l=0.13u
X175 VDD 3bit_freq_divider_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK a_51631_22774# VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0.34p ps=2.68u w=1u l=0.13u
X176 VSS vco_wob_0.vctl a_53086_40850# VSS sg13_lv_nmos ad=0.102p pd=1.28u as=65.99999f ps=0.74u w=0.3u l=0.13u
X177 a_59800_40852# vco_wob_0.vctl VSS VSS sg13_lv_nmos ad=65.99999f pd=0.74u as=0.102p ps=1.28u w=0.3u l=0.13u
X178 VSS a_56887_49467# VSS VSS sg13_lv_nmos ad=95f pd=0.88u as=0 ps=0 w=0.5u l=0.65u
X179 a_53085_40283# a_53022_43738# VDD VDD sg13_lv_pmos ad=59f pd=0.74u as=0.104p ps=1.34u w=0.2u l=0.13u
X180 a_62654_23727# a_61887_24046# a_62270_24055# VSS sg13_lv_nmos ad=0.2017p pd=1.48u as=0.19397p ps=1.29u w=0.64u l=0.13u
X181 3bit_freq_divider_0.EN nEN VDD VDD sg13_lv_pmos ad=0.392p pd=2.94u as=0.392p ps=2.94u w=1.12u l=0.13u
X182 VDD a_58734_56203# a_58734_56203# VDD sg13_lv_pmos ad=0.17p pd=1.68u as=0.17p ps=1.68u w=0.5u l=0.15u
X183 VDD a_64383_23706# a_64817_23685# VDD sg13_lv_pmos ad=79.8f pd=0.8u as=43.05f ps=0.625u w=0.42u l=0.13u
X184 VDD 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.Q a_54472_24641# VDD sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X185 VSS 3bit_freq_divider_0.sg13g2_nand2_1_0.Y 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.sg13g2_dfrbp_1_0.CLK VSS sg13_lv_nmos ad=0.259p pd=2.18u as=0.259p ps=2.18u w=0.74u l=0.13u
X186 a_55862_56737# VDD rhigh l=12u w=1u
X187 VDD a_46817_27899# a_45658_27900# VDD sg13_lv_pmos ad=0.1224p pd=1.4u as=68.39999f ps=0.74u w=0.36u l=0.15u
X188 3bit_freq_divider_1.sg13g2_or3_1_0.B Y1 a_63520_23244# VSS sg13_lv_nmos ad=0.1628p pd=1.18u as=88.8f ps=0.98u w=0.74u l=0.13u
X189 VSS charge_pump_0.vout VSS VSS sg13_lv_nmos ad=0.285p pd=1.88u as=0 ps=0 w=1.5u l=0.65u
X190 a_54489_40413# a_55831_40413# a_55769_40283# VDD sg13_lv_pmos ad=0.1106p pd=0.945u as=0.11p ps=0.94u w=0.5u l=0.13u
X191 a_57084_43159# a_55836_43159# a_57178_43159# VDD sg13_lv_pmos ad=0.17p pd=1.68u as=0.11p ps=0.94u w=0.5u l=0.13u
X192 a_63223_24642# 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.Q VDD VDD sg13_lv_pmos ad=0.1225p pd=1.245u as=0.36p ps=2.72u w=1u l=0.13u
X193 3bit_freq_divider_0.CLK_IN a_57178_43159# a_58426_43159# VDD sg13_lv_pmos ad=0.11p pd=0.94u as=0.11p ps=0.94u w=0.5u l=0.13u
X194 a_58515_40413# 3bit_freq_divider_0.CLK_IN a_59800_40852# VSS sg13_lv_nmos ad=0.11p pd=0.94u as=0.17p ps=1.68u w=0.5u l=0.13u
X195 VDD a_62654_20215# a_62900_20179# VDD sg13_lv_pmos ad=0.2163p pd=1.55u as=79.8f ps=0.8u w=0.42u l=0.13u
X196 a_53086_40850# a_53147_40413# a_52944_43077# VSS sg13_lv_nmos ad=0.17p pd=1.68u as=0.11p ps=0.94u w=0.5u l=0.13u
X197 a_64424_22294# 3bit_freq_divider_1.dff_nclk_0.D a_64424_22200# VSS sg13_lv_nmos ad=50.4f pd=0.66u as=0.1428p ps=1.52u w=0.42u l=0.13u
X198 a_61488_23732# 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.D a_61394_23732# VSS sg13_lv_nmos ad=50.4f pd=0.66u as=0.1428p ps=1.52u w=0.42u l=0.13u
X199 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 3bit_freq_divider_1.sg13g2_nand2_1_0.Y VSS VSS sg13_lv_nmos ad=0.259p pd=2.18u as=0.259p ps=2.18u w=0.74u l=0.13u
X200 a_61061_21478# 3bit_freq_divider_1.freq_div_cell_0.Cout a_60967_21478# VSS sg13_lv_nmos ad=0.1216p pd=1.02u as=0.2176p ps=1.96u w=0.64u l=0.13u
X201 VSS 3bit_freq_divider_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK a_51631_22774# VSS sg13_lv_nmos ad=0.1544p pd=1.235u as=0.2516p ps=2.16u w=0.74u l=0.13u
X202 a_62221_20605# a_61691_20534# a_62119_20605# VDD sg13_lv_pmos ad=51.45f pd=0.665u as=79.8f ps=0.8u w=0.42u l=0.13u
X203 VDD a_53022_43738# a_54427_40283# VDD sg13_lv_pmos ad=0.104p pd=1.34u as=59.75f ps=0.745u w=0.2u l=0.13u
X204 VSS a_53968_22190# a_53899_22244# VSS sg13_lv_nmos ad=0.1825p pd=1.325u as=0.19397p ps=1.29u w=0.64u l=0.13u
X205 VSS charge_pump_0.vout VSS VSS sg13_lv_nmos ad=0.285p pd=1.88u as=0 ps=0 w=1.5u l=0.65u
X206 3bit_freq_divider_1.sg13g2_nand2_1_0.Y 3bit_freq_divider_0.CLK_IN a_60531_21028# VSS sg13_lv_nmos ad=0.2516p pd=2.16u as=66.6f ps=0.92u w=0.74u l=0.13u
X207 VSS a_55345_21385# 3bit_freq_divider_0.freq_div_cell_1.Cout VSS sg13_lv_nmos ad=0.1331p pd=1.12u as=0.2516p ps=2.16u w=0.74u l=0.13u
X208 a_59097_54704# 3bit_freq_divider_0.EN VSS VSS sg13_lv_nmos ad=0.17p pd=1.68u as=0.17p ps=1.68u w=0.5u l=0.15u
X209 a_52114_22293# 3bit_freq_divider_0.dff_nclk_0.D a_51684_22284# VSS sg13_lv_nmos ad=50.4f pd=0.66u as=0.1428p ps=1.52u w=0.42u l=0.13u
X210 a_51693_23075# a_51693_23426# VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0.34p ps=2.68u w=1u l=0.13u
X211 VDD a_64383_23889# a_64383_23706# VDD sg13_lv_pmos ad=0.2163p pd=1.55u as=79.8f ps=0.8u w=0.42u l=0.13u
X212 a_61061_24990# 3bit_freq_divider_1.sg13g2_tiehi_1.L_HI a_60967_24990# VSS sg13_lv_nmos ad=0.1216p pd=1.02u as=0.2176p ps=1.96u w=0.64u l=0.13u
X213 a_58515_40413# VSS cap_cmim l=6.99u w=6.99u
X214 a_54472_21129# 3bit_freq_divider_0.freq_div_cell_0.Cout VDD VDD sg13_lv_pmos ad=0.3808p pd=2.92u as=0.2128p ps=1.5u w=1.12u l=0.13u
X215 a_61887_22290# a_61691_22290# VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0.19p ps=1.38u w=1u l=0.13u
X216 VDD a_53022_43738# a_53058_43159# VDD sg13_lv_pmos ad=0.104p pd=1.34u as=59f ps=0.74u w=0.2u l=0.13u
X217 a_61878_24642# 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.Q VDD VDD sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X218 VSS 3bit_freq_divider_1.dff_nclk_0.nCLK a_61488_21976# VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=50.4f ps=0.66u w=0.42u l=0.13u
X219 a_54400_43159# a_53022_43738# VDD VDD sg13_lv_pmos ad=59f pd=0.74u as=59f ps=0.74u w=0.2u l=0.13u
X220 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.Q a_63463_20216# VSS VSS sg13_lv_nmos ad=0.2516p pd=2.16u as=0.14505p ps=1.15u w=0.74u l=0.13u
X221 a_54434_23148# 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.Q VSS VSS sg13_lv_nmos ad=0.17462p pd=1.185u as=0.15245p ps=1.17u w=0.55u l=0.13u
X222 VDD a_53022_43738# a_55769_40283# VDD sg13_lv_pmos ad=0.104p pd=1.34u as=59.75f ps=0.745u w=0.2u l=0.13u
X223 3bit_freq_divider_0.dff_nclk_0.D a_51648_24041# VDD VDD sg13_lv_pmos ad=0.7616p pd=3.6u as=0.2163p ps=1.55u w=1.12u l=0.13u
X224 3bit_freq_divider_1.freq_div_cell_0.Cout a_60967_23234# VSS VSS sg13_lv_nmos ad=0.2516p pd=2.16u as=0.1331p ps=1.12u w=0.74u l=0.13u
X225 VSS a_56887_49467# VSS VSS sg13_lv_nmos ad=95f pd=0.88u as=0 ps=0 w=0.5u l=0.65u
X226 a_54472_24641# 3bit_freq_divider_0.sg13g2_tiehi_1.L_HI VDD VDD sg13_lv_pmos ad=0.3808p pd=2.92u as=0.2128p ps=1.5u w=1.12u l=0.13u
X227 a_55485_24989# 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.Q VSS VSS sg13_lv_nmos ad=0.1216p pd=1.02u as=0.1331p ps=1.12u w=0.64u l=0.13u
X228 PFD_0.VCO_CLK a_51648_24438# VSS VSS sg13_lv_nmos ad=0.2516p pd=2.16u as=0.14505p ps=1.15u w=0.74u l=0.13u
X229 a_62900_21935# 3bit_freq_divider_1.dff_nclk_0.nCLK VDD VDD sg13_lv_pmos ad=79.8f pd=0.8u as=79.8f ps=0.8u w=0.42u l=0.13u
X230 a_53774_21934# 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0.19p ps=1.38u w=1u l=0.13u
X231 a_55742_43159# a_53022_43738# VDD VDD sg13_lv_pmos ad=59f pd=0.74u as=59f ps=0.74u w=0.2u l=0.13u
X232 a_53899_22244# a_53738_22270# a_53065_21935# VSS sg13_lv_nmos ad=0.19397p pd=1.29u as=0.2017p ps=1.48u w=0.64u l=0.13u
X233 a_64383_23889# a_64383_23628# a_64419_23326# VDD sg13_lv_pmos ad=0.17695p pd=1.56u as=0.19p ps=1.38u w=1u l=0.13u
X234 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.nQ a_62654_23727# VSS VSS sg13_lv_nmos ad=0.2775p pd=2.23u as=0.2516p ps=2.16u w=0.74u l=0.13u
X235 3bit_freq_divider_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 3bit_freq_divider_0.dff_nclk_0.nCLK VDD VDD sg13_lv_pmos ad=0.392p pd=2.94u as=0.392p ps=2.94u w=1.12u l=0.13u
X236 a_58426_43159# a_53022_43738# VDD VDD sg13_lv_pmos ad=59.75f pd=0.745u as=0.104p ps=1.34u w=0.2u l=0.13u
X237 VSS 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.Q a_53054_23243# VSS sg13_lv_nmos ad=0.15245p pd=1.17u as=88.8f ps=0.98u w=0.74u l=0.13u
X238 VSS Y2 a_63255_21488# VSS sg13_lv_nmos ad=0.15245p pd=1.17u as=0.17462p ps=1.185u w=0.55u l=0.13u
X239 VSS a_56887_49467# VSS VSS sg13_lv_nmos ad=95f pd=0.88u as=0 ps=0 w=0.5u l=0.65u
X240 a_52950_20401# a_53065_20179# VDD VDD sg13_lv_pmos ad=0.2856p pd=2.36u as=0.2016p ps=1.5u w=0.84u l=0.13u
X241 a_62119_20605# 3bit_freq_divider_1.dff_nclk_0.nCLK VDD VDD sg13_lv_pmos ad=0.1533p pd=1.57u as=0.11785p ps=1.025u w=0.42u l=0.13u
X242 a_60531_21028# 3bit_freq_divider_0.EN VSS VSS sg13_lv_nmos ad=66.6f pd=0.92u as=0.2516p ps=2.16u w=0.74u l=0.13u
X243 VDD a_52950_20401# 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.Q VDD sg13_lv_pmos ad=0.2016p pd=1.5u as=0.3808p ps=2.92u w=1.12u l=0.13u
X244 a_47777_29803# a_46749_30782# VDD VDD sg13_lv_pmos ad=0.1224p pd=1.4u as=68.39999f ps=0.74u w=0.36u l=0.15u
X245 VSS a_52950_23913# 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.Q VSS sg13_lv_nmos ad=0.14505p pd=1.15u as=0.2516p ps=2.16u w=0.74u l=0.13u
X246 a_51693_23075# a_51693_23426# VSS VSS sg13_lv_nmos ad=0.19397p pd=1.29u as=0.1825p ps=1.325u w=0.64u l=0.13u
X247 VDD 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.sg13g2_dfrbp_1_0.CLK a_61691_24046# VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0.34p ps=2.68u w=1u l=0.13u
X248 a_54602_24999# 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.Q 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.D VSS sg13_lv_nmos ad=88.8f pd=0.98u as=0.1628p ps=1.18u w=0.74u l=0.13u
X249 a_53065_21935# a_53738_22270# a_53702_22368# VDD sg13_lv_pmos ad=0.17695p pd=1.56u as=43.05f ps=0.625u w=0.42u l=0.13u
X250 VSS vco_wob_0.vctl a_53285_42591# VSS sg13_lv_nmos ad=0.102p pd=1.28u as=65.99999f ps=0.74u w=0.3u l=0.13u
X251 VDD a_62654_20215# a_63463_20216# VDD sg13_lv_pmos ad=0.2016p pd=1.5u as=0.2856p ps=2.36u w=0.84u l=0.13u
X252 a_53285_42591# a_52944_43077# a_53152_43159# VSS sg13_lv_nmos ad=0.17p pd=1.68u as=0.11p ps=0.94u w=0.5u l=0.13u
X253 VDD 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.Q a_60967_23234# VDD sg13_lv_pmos ad=0.1918p pd=1.5u as=0.1596p ps=1.22u w=0.84u l=0.13u
X254 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.D a_61707_25000# a_61878_24642# VDD sg13_lv_pmos ad=0.3808p pd=2.92u as=0.2128p ps=1.5u w=1.12u l=0.13u
X255 3bit_freq_divider_1.freq_div_cell_1.Cout a_60967_21478# VDD VDD sg13_lv_pmos ad=0.3808p pd=2.92u as=0.1918p ps=1.5u w=1.12u l=0.13u
X256 a_54842_49733# a_54357_49278# charge_pump_0.vout VDD sg13_lv_pmos ad=55.5f pd=0.74u as=0.1005p ps=1.34u w=0.15u l=0.13u
X257 a_54494_43159# VSS cap_cmim l=6.99u w=6.99u
X258 a_61707_25000# 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.Q a_61675_24642# VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0.1225p ps=1.245u w=1u l=0.13u
X259 a_61394_20220# 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.D VDD VDD sg13_lv_pmos ad=79.8f pd=0.8u as=0.1428p ps=1.52u w=0.42u l=0.13u
X260 VDD 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.D a_54504_22015# VDD sg13_lv_pmos ad=0.1428p pd=1.52u as=79.8f ps=0.8u w=0.42u l=0.13u
X261 a_55345_23141# 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.Q VDD VDD sg13_lv_pmos ad=0.1596p pd=1.22u as=0.1918p ps=1.5u w=0.84u l=0.13u
X262 charge_pump_0.bias_n nEN VSS VSS sg13_lv_nmos ad=0.17p pd=1.68u as=0.17p ps=1.68u w=0.5u l=0.15u
X263 a_53022_43738# a_53022_43738# VDD VDD sg13_lv_pmos ad=59.75f pd=0.745u as=59f ps=0.74u w=0.2u l=0.13u
X264 VSS 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.Q a_61707_25000# VSS sg13_lv_nmos ad=0.15245p pd=1.17u as=0.17462p ps=1.185u w=0.55u l=0.13u
X265 3bit_freq_divider_0.sg13g2_or3_1_0.A a_52886_21392# VSS VSS sg13_lv_nmos ad=0.1628p pd=1.18u as=0.3108p ps=2.32u w=0.74u l=0.13u
X266 VSS charge_pump_0.vout VSS VSS sg13_lv_nmos ad=0.285p pd=1.88u as=0 ps=0 w=1.5u l=0.65u
X267 VSS a_56887_49467# VSS VSS sg13_lv_nmos ad=95f pd=0.88u as=0 ps=0 w=0.5u l=0.65u
X268 a_54427_40283# a_54489_40413# a_53147_40413# VDD sg13_lv_pmos ad=0.17p pd=1.68u as=0.1106p ps=0.945u w=0.5u l=0.13u
X269 a_54252_20259# 3bit_freq_divider_0.dff_nclk_0.nCLK VSS VSS sg13_lv_nmos ad=48.3f pd=0.65u as=0.1825p ps=1.325u w=0.42u l=0.13u
X270 a_54427_40283# a_53022_43738# VDD VDD sg13_lv_pmos ad=59f pd=0.74u as=0.104p ps=1.34u w=0.2u l=0.13u
X271 a_55345_24897# 3bit_freq_divider_0.sg13g2_tiehi_1.L_HI a_55485_24989# VSS sg13_lv_nmos ad=0.2176p pd=1.96u as=0.1216p ps=1.02u w=0.64u l=0.13u
X272 CLK_OUT a_64384_24445# VSS VSS sg13_lv_nmos ad=0.2516p pd=2.16u as=0.14505p ps=1.15u w=0.74u l=0.13u
X273 a_54504_20259# a_53774_20178# a_53968_20434# VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=79.8f ps=0.8u w=0.42u l=0.13u
X274 VSS charge_pump_0.vout VSS VSS sg13_lv_nmos ad=0.285p pd=1.88u as=0 ps=0 w=1.5u l=0.65u
X275 VSS a_51685_23725# a_52119_23653# VSS sg13_lv_nmos ad=90.3f pd=0.85u as=54.6f ps=0.68u w=0.42u l=0.13u
X276 VDD 3bit_freq_divider_1.freq_div_cell_0.Cout a_61878_21130# VDD sg13_lv_pmos ad=0.2128p pd=1.5u as=0.3808p ps=2.92u w=1.12u l=0.13u
X277 a_52950_22157# a_53065_21935# VSS VSS sg13_lv_nmos ad=0.187p pd=1.78u as=0.14505p ps=1.15u w=0.55u l=0.13u
X278 a_55969_42591# vco_wob_0.vctl VSS VSS sg13_lv_nmos ad=65.99999f pd=0.74u as=0.102p ps=1.28u w=0.3u l=0.13u
X279 a_55836_43159# a_54494_43159# a_55969_42591# VSS sg13_lv_nmos ad=0.11p pd=0.94u as=0.17p ps=1.68u w=0.5u l=0.13u
X280 a_55770_40850# vco_wob_0.vctl VSS VSS sg13_lv_nmos ad=65.99999f pd=0.74u as=0.102p ps=1.28u w=0.3u l=0.13u
X281 a_62654_23727# a_61691_24046# a_62270_24055# VDD sg13_lv_pmos ad=0.17695p pd=1.56u as=0.19p ps=1.38u w=1u l=0.13u
X282 a_64714_21414# 3bit_freq_divider_1.sg13g2_or3_1_0.B a_64714_21300# VDD sg13_lv_pmos ad=0.1275p pd=1.255u as=0.22p ps=1.44u w=1u l=0.13u
X283 VDD a_51648_24041# a_51648_24438# VDD sg13_lv_pmos ad=0.2016p pd=1.5u as=0.2856p ps=2.36u w=0.84u l=0.13u
X284 VSS a_56887_49467# VSS VSS sg13_lv_nmos ad=95f pd=0.88u as=0 ps=0 w=0.5u l=0.65u
X285 a_55831_40413# VSS cap_cmim l=6.99u w=6.99u
X286 a_52924_21129# 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.Q VDD VDD sg13_lv_pmos ad=0.3808p pd=2.92u as=0.2128p ps=1.5u w=1.12u l=0.13u
X287 VSS a_56887_49467# VSS VSS sg13_lv_nmos ad=95f pd=0.88u as=0 ps=0 w=0.5u l=0.65u
X288 a_55769_40283# a_55831_40413# a_54489_40413# VDD sg13_lv_pmos ad=0.17p pd=1.68u as=0.1106p ps=0.945u w=0.5u l=0.13u
X289 VSS a_62654_21971# a_63463_21972# VSS sg13_lv_nmos ad=0.14505p pd=1.15u as=0.187p ps=1.78u w=0.55u l=0.13u
X290 a_54252_23771# 3bit_freq_divider_0.dff_nclk_0.nCLK VSS VSS sg13_lv_nmos ad=48.3f pd=0.65u as=0.1825p ps=1.325u w=0.42u l=0.13u
X291 VDD a_45658_27900# PFD_0.DOWN VDD sg13_lv_pmos ad=0.1088p pd=1.32u as=60.8f ps=0.7u w=0.32u l=0.15u
X292 3bit_freq_divider_1.dff_nclk_0.D a_64383_23889# VDD VDD sg13_lv_pmos ad=0.7616p pd=3.6u as=0.2163p ps=1.55u w=1.12u l=0.13u
X293 a_45658_27900# a_46817_27899# VDD VDD sg13_lv_pmos ad=68.39999f pd=0.74u as=0.1224p ps=1.4u w=0.36u l=0.15u
X294 VSS 3bit_freq_divider_0.dff_nclk_0.nCLK a_53539_21970# VSS sg13_lv_nmos ad=90.3f pd=0.85u as=47.25f ps=0.645u w=0.42u l=0.13u
X295 a_53539_21970# a_53065_21935# a_53445_21970# VSS sg13_lv_nmos ad=47.25f pd=0.645u as=0.1428p ps=1.52u w=0.42u l=0.13u
X296 VDD 3bit_freq_divider_0.dff_nclk_0.nCLK a_53968_22190# VDD sg13_lv_pmos ad=0.11785p pd=1.025u as=0.1533p ps=1.57u w=0.42u l=0.13u
X297 a_54504_23771# a_53774_23690# a_53968_23946# VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=79.8f ps=0.8u w=0.42u l=0.13u
X298 VSS a_53968_23946# a_53899_24000# VSS sg13_lv_nmos ad=0.1825p pd=1.325u as=0.19397p ps=1.29u w=0.64u l=0.13u
X299 a_52924_22885# a_52886_23148# 3bit_freq_divider_0.sg13g2_or3_1_0.B VDD sg13_lv_pmos ad=0.2128p pd=1.5u as=0.3808p ps=2.92u w=1.12u l=0.13u
X300 a_52886_23148# X1 VSS VSS sg13_lv_nmos ad=0.17462p pd=1.185u as=0.15245p ps=1.17u w=0.55u l=0.13u
X301 a_58453_40283# a_58515_40413# a_57173_40413# VDD sg13_lv_pmos ad=0.11p pd=0.94u as=0.11p ps=0.94u w=0.5u l=0.13u
X302 a_63520_21488# 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.Q VSS VSS sg13_lv_nmos ad=88.8f pd=0.98u as=0.15245p ps=1.17u w=0.74u l=0.13u
X303 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.nQ a_62654_23727# VDD VDD sg13_lv_pmos ad=0.7616p pd=3.6u as=0.2163p ps=1.55u w=1.12u l=0.13u
X304 a_54427_40283# a_53022_43738# VDD VDD sg13_lv_pmos ad=59.75f pd=0.745u as=59f ps=0.74u w=0.2u l=0.13u
X305 a_64731_24890# a_64398_24796# 3bit_freq_divider_1.dff_nclk_0.nRST VDD sg13_lv_pmos ad=0.4657p pd=2.54u as=0.3927p ps=2.99u w=1.155u l=0.13u
X306 a_61707_21488# 3bit_freq_divider_1.freq_div_cell_0.Cout VSS VSS sg13_lv_nmos ad=0.17462p pd=1.185u as=0.374p ps=2.46u w=0.55u l=0.13u
X307 VDD a_53968_22190# a_53899_22244# VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0.19p ps=1.38u w=1u l=0.13u
X308 VSS a_56887_49467# VSS VSS sg13_lv_nmos ad=95f pd=0.88u as=0 ps=0 w=0.5u l=0.65u
X309 a_52924_24641# 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.Q VDD VDD sg13_lv_pmos ad=0.3808p pd=2.92u as=0.2128p ps=1.5u w=1.12u l=0.13u
X310 VSS a_56887_49467# VSS VSS sg13_lv_nmos ad=95f pd=0.88u as=0 ps=0 w=0.5u l=0.65u
X311 a_54489_40413# a_55831_40413# a_55770_40850# VSS sg13_lv_nmos ad=0.11p pd=0.94u as=0.17p ps=1.68u w=0.5u l=0.13u
X312 VDD a_52950_23913# 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.Q VDD sg13_lv_pmos ad=0.2016p pd=1.5u as=0.3808p ps=2.92u w=1.12u l=0.13u
X313 a_61887_24046# a_61691_24046# VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0.19p ps=1.38u w=1u l=0.13u
X314 charge_pump_0.vout vco_wob_0.vctl rhigh l=0.96u w=0.6u
X315 VDD a_53065_21935# 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.nQ VDD sg13_lv_pmos ad=0.2163p pd=1.55u as=0.7616p ps=3.6u w=1.12u l=0.13u
X316 a_53152_43159# a_52944_43077# a_53058_43159# VDD sg13_lv_pmos ad=0.11p pd=0.94u as=0.11p ps=0.94u w=0.5u l=0.13u
X317 VDD a_51685_23725# a_51721_23684# VDD sg13_lv_pmos ad=79.8f pd=0.8u as=43.05f ps=0.625u w=0.42u l=0.13u
X318 VDD a_53774_23690# a_53738_24026# VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0.34p ps=2.68u w=1u l=0.13u
X319 a_55836_43159# a_54494_43159# a_55742_43159# VDD sg13_lv_pmos ad=0.1106p pd=0.945u as=0.17p ps=1.68u w=0.5u l=0.13u
X320 a_55769_40283# a_53022_43738# VDD VDD sg13_lv_pmos ad=59.75f pd=0.745u as=59f ps=0.74u w=0.2u l=0.13u
X321 a_56013_24979# a_56137_24678# a_56038_24617# VDD sg13_lv_pmos ad=0.2442p pd=2.06u as=0.4657p ps=2.54u w=0.66u l=0.13u
X322 VDD 3bit_freq_divider_0.freq_div_cell_0.Cin a_55345_23141# VDD sg13_lv_pmos ad=0.2856p pd=2.36u as=0.1596p ps=1.22u w=0.84u l=0.13u
X323 VSS a_56887_49467# VSS VSS sg13_lv_nmos ad=95f pd=0.88u as=0 ps=0 w=0.5u l=0.65u
X324 a_48909_28913# CLK_IN VSS VSS sg13_lv_nmos ad=0.1224p pd=1.4u as=0.1224p ps=1.4u w=0.36u l=0.15u
X325 a_64464_23052# a_64383_23434# a_64383_23300# VSS sg13_lv_nmos ad=54.6f pd=0.68u as=79.8f ps=0.8u w=0.42u l=0.13u
X326 a_56055_21027# 3bit_freq_divider_0.CLK_IN 3bit_freq_divider_0.sg13g2_nand2_1_0.Y VSS sg13_lv_nmos ad=66.6f pd=0.92u as=0.2516p ps=2.16u w=0.74u l=0.13u
X327 VSS a_56887_49467# VSS VSS sg13_lv_nmos ad=95f pd=0.88u as=0 ps=0 w=0.5u l=0.65u
X328 a_61972_25000# 3bit_freq_divider_1.sg13g2_tiehi_1.L_HI VSS VSS sg13_lv_nmos ad=88.8f pd=0.98u as=0.15245p ps=1.17u w=0.74u l=0.13u
X329 a_63255_21488# Y2 a_63223_21130# VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0.1225p ps=1.245u w=1u l=0.13u
X330 a_51648_21103# 3bit_freq_divider_0.sg13g2_or3_1_0.C VSS VSS sg13_lv_nmos ad=0.187p pd=1.78u as=0.1045p ps=0.93u w=0.55u l=0.13u
X331 a_53899_24000# a_53738_24026# a_53065_23691# VSS sg13_lv_nmos ad=0.19397p pd=1.29u as=0.2017p ps=1.48u w=0.64u l=0.13u
X332 VSS 3bit_freq_divider_0.freq_div_cell_0.Cin a_54434_23148# VSS sg13_lv_nmos ad=0.374p pd=2.46u as=0.17462p ps=1.185u w=0.55u l=0.13u
X333 charge_pump_0.vout PFD_0.DOWN a_54747_49259# VSS sg13_lv_nmos ad=0.408p pd=3.08u as=0.207p ps=1.545u w=1.2u l=0.13u
X334 a_52119_23843# 3bit_freq_divider_0.dff_nclk_0.nRST VSS VSS sg13_lv_nmos ad=47.25f pd=0.645u as=90.3f ps=0.85u w=0.42u l=0.13u
X335 PFD_0.UP a_47777_29803# VDD VDD sg13_lv_pmos ad=0.1088p pd=1.32u as=60.8f ps=0.7u w=0.32u l=0.15u
X336 a_53054_24999# X0 3bit_freq_divider_0.sg13g2_or3_1_0.C VSS sg13_lv_nmos ad=88.8f pd=0.98u as=0.1628p ps=1.18u w=0.74u l=0.13u
X337 VSS charge_pump_0.vout VSS VSS sg13_lv_nmos ad=0.285p pd=1.88u as=0 ps=0 w=1.5u l=0.65u
X338 a_57178_43159# a_55836_43159# a_57084_43159# VDD sg13_lv_pmos ad=0.1106p pd=0.945u as=0.17p ps=1.68u w=0.5u l=0.13u
X339 VDD a_55345_21385# 3bit_freq_divider_0.freq_div_cell_1.Cout VDD sg13_lv_pmos ad=0.1918p pd=1.5u as=0.3808p ps=2.92u w=1.12u l=0.13u
X340 VDD 3bit_freq_divider_1.dff_nclk_0.nCLK a_61394_23732# VDD sg13_lv_pmos ad=0.1428p pd=1.52u as=79.8f ps=0.8u w=0.42u l=0.13u
X341 VSS a_56887_49467# VSS VSS sg13_lv_nmos ad=95f pd=0.88u as=0 ps=0 w=0.5u l=0.65u
X342 a_57084_43159# a_53022_43738# VDD VDD sg13_lv_pmos ad=59f pd=0.74u as=59f ps=0.74u w=0.2u l=0.13u
X343 a_53065_21935# a_53774_21934# a_53722_21970# VSS sg13_lv_nmos ad=0.2017p pd=1.48u as=54.6f ps=0.68u w=0.42u l=0.13u
X344 a_53968_22190# a_53774_21934# a_54352_22360# VDD sg13_lv_pmos ad=79.8f pd=0.8u as=51.45f ps=0.665u w=0.42u l=0.13u
X345 a_53702_20612# a_53445_20214# VDD VDD sg13_lv_pmos ad=43.05f pd=0.625u as=79.8f ps=0.8u w=0.42u l=0.13u
X346 VDD a_53022_43738# a_58426_43159# VDD sg13_lv_pmos ad=59f pd=0.74u as=59.75f ps=0.745u w=0.2u l=0.13u
X347 VSS vco_wob_0.vctl a_59800_40852# VSS sg13_lv_nmos ad=0.102p pd=1.28u as=65.99999f ps=0.74u w=0.3u l=0.13u
X348 a_59799_40285# a_53022_43738# VDD VDD sg13_lv_pmos ad=59f pd=0.74u as=0.104p ps=1.34u w=0.2u l=0.13u
X349 a_60967_24990# 3bit_freq_divider_1.sg13g2_tiehi_1.L_HI VDD VDD sg13_lv_pmos ad=0.1596p pd=1.22u as=0.2856p ps=2.36u w=0.84u l=0.13u
X350 VDD a_53022_43738# a_53085_40283# VDD sg13_lv_pmos ad=59f pd=0.74u as=59f ps=0.74u w=0.2u l=0.13u
X351 a_53722_21970# a_53445_21970# VSS VSS sg13_lv_nmos ad=54.6f pd=0.68u as=90.3f ps=0.85u w=0.42u l=0.13u
X352 VSS charge_pump_0.vout VSS VSS sg13_lv_nmos ad=0.285p pd=1.88u as=0 ps=0 w=1.5u l=0.65u
X353 VSS vco_wob_0.vctl a_54428_40850# VSS sg13_lv_nmos ad=0.102p pd=1.28u as=65.99999f ps=0.74u w=0.3u l=0.13u
X354 VSS charge_pump_0.vout VSS VSS sg13_lv_nmos ad=0.285p pd=1.88u as=0 ps=0 w=1.5u l=0.65u
X355 VSS 3bit_freq_divider_1.dff_nclk_0.nCLK a_62324_23772# VSS sg13_lv_nmos ad=0.1825p pd=1.325u as=48.3f ps=0.65u w=0.42u l=0.13u
X356 VDD a_55345_24897# 3bit_freq_divider_0.freq_div_cell_0.Cin VDD sg13_lv_pmos ad=0.1918p pd=1.5u as=0.3808p ps=2.92u w=1.12u l=0.13u
X357 VSS a_63255_23244# 3bit_freq_divider_1.sg13g2_or3_1_0.B VSS sg13_lv_nmos ad=0.3108p pd=2.32u as=0.1628p ps=1.18u w=0.74u l=0.13u
X358 a_61675_24642# 3bit_freq_divider_1.sg13g2_tiehi_1.L_HI VDD VDD sg13_lv_pmos ad=0.1225p pd=1.245u as=0.36p ps=2.72u w=1u l=0.13u
X359 a_53058_43159# a_53022_43738# VDD VDD sg13_lv_pmos ad=59.75f pd=0.745u as=0.104p ps=1.34u w=0.2u l=0.13u
X360 VDD 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.Q a_63426_22886# VDD sg13_lv_pmos ad=0.2128p pd=1.5u as=0.3808p ps=2.92u w=1.12u l=0.13u
X361 3bit_freq_divider_0.sg13g2_nand2_1_0.Y 3bit_freq_divider_0.CLK_IN VDD VDD sg13_lv_pmos ad=0.2128p pd=1.5u as=0.3808p ps=2.92u w=1.12u l=0.13u
X362 a_53968_22190# a_53738_22270# a_54324_22015# VSS sg13_lv_nmos ad=79.8f pd=0.8u as=54.6f ps=0.68u w=0.42u l=0.13u
X363 a_63426_21130# Y2 VDD VDD sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X364 a_57173_40413# VSS cap_cmim l=6.99u w=6.99u
X365 a_61394_21976# 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.D VDD VDD sg13_lv_pmos ad=79.8f pd=0.8u as=0.1428p ps=1.52u w=0.42u l=0.13u
X366 VSS charge_pump_0.vout VSS VSS sg13_lv_nmos ad=0.285p pd=1.88u as=0 ps=0 w=1.5u l=0.65u
X367 a_54324_22015# a_53899_22244# a_54252_22015# VSS sg13_lv_nmos ad=54.6f pd=0.68u as=48.3f ps=0.65u w=0.42u l=0.13u
X368 a_59800_40852# 3bit_freq_divider_0.CLK_IN a_58515_40413# VSS sg13_lv_nmos ad=0.17p pd=1.68u as=0.11p ps=0.94u w=0.5u l=0.13u
X369 a_58734_56203# a_58536_54976# a_58536_54976# VDD sg13_lv_pmos ad=0.17p pd=1.68u as=0.17p ps=1.68u w=0.5u l=0.15u
X370 a_54428_40850# a_54489_40413# a_53147_40413# VSS sg13_lv_nmos ad=0.17p pd=1.68u as=0.11p ps=0.94u w=0.5u l=0.13u
X371 a_52950_23913# a_53065_23691# VSS VSS sg13_lv_nmos ad=0.187p pd=1.78u as=0.14505p ps=1.15u w=0.55u l=0.13u
X372 a_64383_23300# a_64383_23434# a_64424_22200# VDD sg13_lv_pmos ad=79.8f pd=0.8u as=0.1428p ps=1.52u w=0.42u l=0.13u
X373 VSS 3bit_freq_divider_1.sg13g2_or3_1_0.B a_64384_21091# VSS sg13_lv_nmos ad=0.1045p pd=0.93u as=0.198p ps=1.27u w=0.55u l=0.13u
X374 VSS 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.Q a_52886_24904# VSS sg13_lv_nmos ad=0.374p pd=2.46u as=0.17462p ps=1.185u w=0.55u l=0.13u
X375 VDD 3bit_freq_divider_0.dff_nclk_0.nRST a_51684_22284# VDD sg13_lv_pmos ad=0.1428p pd=1.52u as=79.8f ps=0.8u w=0.42u l=0.13u
X376 VDD charge_pump_0.bias_p charge_pump_0.bias_p VDD sg13_lv_pmos ad=0.68p pd=4.68u as=0.68p ps=4.68u w=2u l=1u
X377 a_64459_24995# a_64459_24995# a_64338_24910# VSS sg13_lv_nmos ad=0.102p pd=1.28u as=0.2307p ps=1.615u w=0.3u l=0.13u
X378 VDD 3bit_freq_divider_0.dff_nclk_0.nCLK a_53445_21970# VDD sg13_lv_pmos ad=79.8f pd=0.8u as=79.8f ps=0.8u w=0.42u l=0.13u
X379 VDD PFD_0.UP a_54357_49278# VDD sg13_lv_pmos ad=0.102p pd=1.28u as=0.102p ps=1.28u w=0.3u l=0.13u
X380 VSS a_62654_23727# a_63463_23728# VSS sg13_lv_nmos ad=0.14505p pd=1.15u as=0.187p ps=1.78u w=0.55u l=0.13u
X381 VSS charge_pump_0.vout VSS VSS sg13_lv_nmos ad=0.285p pd=1.88u as=0 ps=0 w=1.5u l=0.65u
X382 a_53899_24000# a_53774_23690# a_53065_23691# VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0.17695p ps=1.56u w=1u l=0.13u
X383 VDD 3bit_freq_divider_0.dff_nclk_0.nCLK a_53968_23946# VDD sg13_lv_pmos ad=0.11785p pd=1.025u as=0.1533p ps=1.57u w=0.42u l=0.13u
X384 a_53539_23726# a_53065_23691# a_53445_23726# VSS sg13_lv_nmos ad=47.25f pd=0.645u as=0.1428p ps=1.52u w=0.42u l=0.13u
X385 VSS 3bit_freq_divider_0.dff_nclk_0.nCLK a_53539_23726# VSS sg13_lv_nmos ad=90.3f pd=0.85u as=47.25f ps=0.645u w=0.42u l=0.13u
X386 a_57311_42591# vco_wob_0.vctl VSS VSS sg13_lv_nmos ad=65.99999f pd=0.74u as=0.102p ps=1.28u w=0.3u l=0.13u
X387 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.D 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.Q a_61972_25000# VSS sg13_lv_nmos ad=0.1628p pd=1.18u as=88.8f ps=0.98u w=0.74u l=0.13u
X388 3bit_freq_divider_1.sg13g2_or3_1_0.C a_63255_25000# a_63426_24642# VDD sg13_lv_pmos ad=0.3808p pd=2.92u as=0.2128p ps=1.5u w=1.12u l=0.13u
X389 a_57178_43159# a_55836_43159# a_57311_42591# VSS sg13_lv_nmos ad=0.11p pd=0.94u as=0.17p ps=1.68u w=0.5u l=0.13u
X390 a_45579_29803# CLK_IN a_45451_28860# VSS sg13_lv_nmos ad=0.1224p pd=1.4u as=68.39999f ps=0.74u w=0.36u l=0.15u
X391 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.Q a_63463_21972# VDD VDD sg13_lv_pmos ad=0.3808p pd=2.92u as=0.2016p ps=1.5u w=1.12u l=0.13u
X392 VSS 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.sg13g2_dfrbp_1_0.CLK a_61691_24046# VSS sg13_lv_nmos ad=0.1544p pd=1.235u as=0.2516p ps=2.16u w=0.74u l=0.13u
X393 VDD 3bit_freq_divider_1.dff_nclk_0.nRST a_64424_22200# VDD sg13_lv_pmos ad=0.1428p pd=1.52u as=79.8f ps=0.8u w=0.42u l=0.13u
X394 VDD a_64419_23326# a_64809_23027# VDD sg13_lv_pmos ad=0.11785p pd=1.025u as=51.45f ps=0.665u w=0.42u l=0.13u
X395 a_64338_24910# a_64362_24865# a_64398_24796# VSS sg13_lv_nmos ad=0.2307p pd=1.615u as=0.27427p ps=2.28u w=0.795u l=0.13u
X396 a_62654_20215# a_61887_20534# a_62270_20543# VSS sg13_lv_nmos ad=0.2017p pd=1.48u as=0.19397p ps=1.29u w=0.64u l=0.13u
X397 PFD_0.DOWN a_45658_27900# VDD VDD sg13_lv_pmos ad=60.8f pd=0.7u as=60.8f ps=0.7u w=0.32u l=0.15u
X398 a_54472_22885# a_54434_23148# 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.D VDD sg13_lv_pmos ad=0.2128p pd=1.5u as=0.3808p ps=2.92u w=1.12u l=0.13u
X399 VDD 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.Q a_53350_22885# VDD sg13_lv_pmos ad=0.36p pd=2.72u as=0.1225p ps=1.245u w=1u l=0.13u
X400 VSS 3bit_freq_divider_0.sg13g2_nand2_1_0.Y 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.sg13g2_dfrbp_1_0.CLK VSS sg13_lv_nmos ad=0.259p pd=2.18u as=0.259p ps=2.18u w=0.74u l=0.13u
X401 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 3bit_freq_divider_1.sg13g2_nand2_1_0.Y VDD VDD sg13_lv_pmos ad=0.392p pd=2.94u as=0.392p ps=2.94u w=1.12u l=0.13u
X402 a_51648_24041# a_51684_22692# a_51693_23075# VSS sg13_lv_nmos ad=0.2017p pd=1.48u as=0.19397p ps=1.29u w=0.64u l=0.13u
X403 VDD a_62900_23691# a_62879_24125# VDD sg13_lv_pmos ad=79.8f pd=0.8u as=43.05f ps=0.625u w=0.42u l=0.13u
X404 VSS 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.Q a_61707_21488# VSS sg13_lv_nmos ad=0.15245p pd=1.17u as=0.17462p ps=1.185u w=0.55u l=0.13u
X405 a_45579_29803# CLK_IN a_45451_28860# VSS sg13_lv_nmos ad=68.39999f pd=0.74u as=68.39999f ps=0.74u w=0.36u l=0.15u
X406 VSS 3bit_freq_divider_1.dff_nclk_0.nRST a_64424_22294# VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=50.4f ps=0.66u w=0.42u l=0.13u
X407 a_45579_29803# CLK_IN VDD VDD sg13_lv_pmos ad=0.1088p pd=1.32u as=60.8f ps=0.7u w=0.32u l=0.15u
X408 VSS 3bit_freq_divider_0.sg13g2_tiehi_1.L_HI a_54602_24999# VSS sg13_lv_nmos ad=0.15245p pd=1.17u as=88.8f ps=0.98u w=0.74u l=0.13u
X409 a_63223_21130# 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.Q VDD VDD sg13_lv_pmos ad=0.1225p pd=1.245u as=0.36p ps=2.72u w=1u l=0.13u
X410 a_58515_40413# 3bit_freq_divider_0.CLK_IN a_59799_40285# VDD sg13_lv_pmos ad=0.11p pd=0.94u as=0.17p ps=1.68u w=0.5u l=0.13u
X411 a_53085_40283# a_53147_40413# a_52944_43077# VDD sg13_lv_pmos ad=0.11p pd=0.94u as=0.11p ps=0.94u w=0.5u l=0.13u
X412 a_58515_40413# 3bit_freq_divider_0.CLK_IN a_59799_40285# VDD sg13_lv_pmos ad=0.1106p pd=0.945u as=0.11p ps=0.94u w=0.5u l=0.13u
X413 a_61488_20220# 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.D a_61394_20220# VSS sg13_lv_nmos ad=50.4f pd=0.66u as=0.1428p ps=1.52u w=0.42u l=0.13u
X414 a_62654_20215# a_61691_20534# a_62270_20543# VDD sg13_lv_pmos ad=0.17695p pd=1.56u as=0.19p ps=1.38u w=1u l=0.13u
X415 a_54494_43159# a_53152_43159# a_54400_43159# VDD sg13_lv_pmos ad=0.11p pd=0.94u as=0.11p ps=0.94u w=0.5u l=0.13u
X416 VSS charge_pump_0.vout VSS VSS sg13_lv_nmos ad=0.285p pd=1.88u as=0 ps=0 w=1.5u l=0.65u
X417 a_55742_43159# a_54494_43159# a_55836_43159# VDD sg13_lv_pmos ad=0.11p pd=0.94u as=0.1106p ps=0.945u w=0.5u l=0.13u
X418 a_46817_27899# PFD_0.VCO_CLK a_47954_28913# VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=79.8f ps=0.8u w=0.42u l=0.15u
X419 VSS 3bit_freq_divider_0.dff_nclk_0.nRST a_52114_22293# VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=50.4f ps=0.66u w=0.42u l=0.13u
X420 VSS a_53065_21935# 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.nQ VSS sg13_lv_nmos ad=0.2516p pd=2.16u as=0.2775p ps=2.23u w=0.74u l=0.13u
X421 VDD a_53022_43738# a_58453_40283# VDD sg13_lv_pmos ad=59f pd=0.74u as=59f ps=0.74u w=0.2u l=0.13u
X422 a_54352_22360# a_53899_22244# VDD VDD sg13_lv_pmos ad=51.45f pd=0.665u as=0.11785p ps=1.025u w=0.42u l=0.13u
X423 VSS a_61707_23244# 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.D VSS sg13_lv_nmos ad=0.3108p pd=2.32u as=0.1628p ps=1.18u w=0.74u l=0.13u
X424 a_54357_49278# PFD_0.UP VSS VSS sg13_lv_nmos ad=0.1005p pd=1.34u as=0.1005p ps=1.34u w=0.15u l=0.13u
X425 a_53968_23946# a_53774_23690# a_54352_24116# VDD sg13_lv_pmos ad=79.8f pd=0.8u as=51.45f ps=0.665u w=0.42u l=0.13u
X426 VDD 3bit_freq_divider_0.sg13g2_nand2_1_0.Y 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK VDD sg13_lv_pmos ad=0.392p pd=2.94u as=0.392p ps=2.94u w=1.12u l=0.13u
X427 VSS a_56887_49467# VSS VSS sg13_lv_nmos ad=0.17p pd=1.68u as=0 ps=0 w=0.5u l=0.65u
X428 a_53065_23691# a_53774_23690# a_53722_23726# VSS sg13_lv_nmos ad=0.2017p pd=1.48u as=54.6f ps=0.68u w=0.42u l=0.13u
X429 a_61878_21130# 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.Q VDD VDD sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X430 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.D a_54434_23148# VSS VSS sg13_lv_nmos ad=0.1628p pd=1.18u as=0.3108p ps=2.32u w=0.74u l=0.13u
X431 VDD 3bit_freq_divider_0.EN a_58536_54976# VDD sg13_lv_pmos ad=0.17p pd=1.68u as=0.17p ps=1.68u w=0.5u l=0.15u
X432 a_57084_43159# a_55836_43159# a_57178_43159# VDD sg13_lv_pmos ad=0.11p pd=0.94u as=0.1106p ps=0.945u w=0.5u l=0.13u
X433 VDD 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.sg13g2_dfrbp_1_0.CLK a_61691_20534# VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0.34p ps=2.68u w=1u l=0.13u
X434 a_53722_23726# a_53445_23726# VSS VSS sg13_lv_nmos ad=54.6f pd=0.68u as=90.3f ps=0.85u w=0.42u l=0.13u
X435 a_55086_20219# 3bit_freq_divider_0.dff_nclk_0.nCLK VSS VSS sg13_lv_nmos ad=50.4f pd=0.66u as=0.1428p ps=1.52u w=0.42u l=0.13u
X436 3bit_freq_divider_0.CLK_IN VSS cap_cmim l=6.99u w=6.99u
X437 3bit_freq_divider_0.CLK_IN a_57178_43159# a_58426_43159# VDD sg13_lv_pmos ad=0.1106p pd=0.945u as=0.17p ps=1.68u w=0.5u l=0.13u
X438 PFD_0.UP a_47777_29803# VDD VDD sg13_lv_pmos ad=60.8f pd=0.7u as=0.1088p ps=1.32u w=0.32u l=0.15u
X439 a_62879_22369# a_61887_22290# a_62654_21971# VDD sg13_lv_pmos ad=43.05f pd=0.625u as=0.17695p ps=1.56u w=0.42u l=0.13u
X440 VDD a_47777_29803# PFD_0.UP VDD sg13_lv_pmos ad=60.8f pd=0.7u as=60.8f ps=0.7u w=0.32u l=0.15u
X441 VSS 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.Q a_61061_21478# VSS sg13_lv_nmos ad=0.1331p pd=1.12u as=0.1216p ps=1.02u w=0.64u l=0.13u
X442 a_51600_24907# a_51622_24863# 3bit_freq_divider_0.dff_nclk_0.nRST VDD sg13_lv_pmos ad=0.4657p pd=2.54u as=0.3927p ps=2.99u w=1.155u l=0.13u
X443 VSS 3bit_freq_divider_1.dff_nclk_0.nRST a_64464_23130# VSS sg13_lv_nmos ad=0.1825p pd=1.325u as=48.3f ps=0.65u w=0.42u l=0.13u
X444 VSS a_56887_49467# VSS VSS sg13_lv_nmos ad=0.17p pd=1.68u as=0 ps=0 w=0.5u l=0.65u
X445 VDD a_46749_30782# a_47777_29803# VDD sg13_lv_pmos ad=68.39999f pd=0.74u as=0.1224p ps=1.4u w=0.36u l=0.15u
X446 a_55485_21477# 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.Q VSS VSS sg13_lv_nmos ad=0.1216p pd=1.02u as=0.1331p ps=1.12u w=0.64u l=0.13u
X447 VSS a_56887_49467# VSS VSS sg13_lv_nmos ad=95f pd=0.88u as=0 ps=0 w=0.5u l=0.65u
X448 VSS vco_wob_0.vctl a_55969_42591# VSS sg13_lv_nmos ad=0.102p pd=1.28u as=65.99999f ps=0.74u w=0.3u l=0.13u
X449 a_55969_42591# a_54494_43159# a_55836_43159# VSS sg13_lv_nmos ad=0.17p pd=1.68u as=0.11p ps=0.94u w=0.5u l=0.13u
X450 VSS vco_wob_0.vctl a_55770_40850# VSS sg13_lv_nmos ad=0.102p pd=1.28u as=65.99999f ps=0.74u w=0.3u l=0.13u
X451 a_53022_43738# vco_wob_0.vctl VSS VSS sg13_lv_nmos ad=65.99999f pd=0.74u as=0.102p ps=1.28u w=0.3u l=0.13u
X452 a_55769_40283# a_53022_43738# VDD VDD sg13_lv_pmos ad=59f pd=0.74u as=0.104p ps=1.34u w=0.2u l=0.13u
X453 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.nQ a_62654_20215# VSS VSS sg13_lv_nmos ad=0.2775p pd=2.23u as=0.2516p ps=2.16u w=0.74u l=0.13u
X454 a_55086_23731# 3bit_freq_divider_0.dff_nclk_0.nCLK VSS VSS sg13_lv_nmos ad=50.4f pd=0.66u as=0.1428p ps=1.52u w=0.42u l=0.13u
X455 VSS 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.Q a_61061_24990# VSS sg13_lv_nmos ad=0.1331p pd=1.12u as=0.1216p ps=1.02u w=0.64u l=0.13u
X456 VSS a_64383_23706# a_64419_23654# VSS sg13_lv_nmos ad=90.3f pd=0.85u as=54.6f ps=0.68u w=0.42u l=0.13u
X457 a_61972_21488# 3bit_freq_divider_1.freq_div_cell_0.Cout VSS VSS sg13_lv_nmos ad=88.8f pd=0.98u as=0.15245p ps=1.17u w=0.74u l=0.13u
X458 VDD a_53022_43738# a_53058_43159# VDD sg13_lv_pmos ad=59f pd=0.74u as=59.75f ps=0.745u w=0.2u l=0.13u
X459 VSS vco_wob_0.vctl VSS VSS sg13_lv_nmos ad=0.1005p pd=1.34u as=0 ps=0 w=0.15u l=0.13u
X460 a_54434_24904# 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.Q VSS VSS sg13_lv_nmos ad=0.17462p pd=1.185u as=0.15245p ps=1.17u w=0.55u l=0.13u
X461 a_53445_23726# a_53065_23691# VDD VDD sg13_lv_pmos ad=79.8f pd=0.8u as=0.2163p ps=1.55u w=0.42u l=0.13u
X462 a_54400_43159# a_53022_43738# VDD VDD sg13_lv_pmos ad=59.75f pd=0.745u as=0.104p ps=1.34u w=0.2u l=0.13u
X463 a_51684_22692# a_51631_22774# VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0.19p ps=1.38u w=1u l=0.13u
X464 VSS a_56887_49467# VSS VSS sg13_lv_nmos ad=95f pd=0.88u as=0 ps=0 w=0.5u l=0.65u
X465 a_57111_40283# a_57173_40413# a_55831_40413# VDD sg13_lv_pmos ad=0.17p pd=1.68u as=0.1106p ps=0.945u w=0.5u l=0.13u
X466 a_63255_25000# 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.Q VSS VSS sg13_lv_nmos ad=0.17462p pd=1.185u as=0.374p ps=2.46u w=0.55u l=0.13u
X467 charge_pump_0.bias_p a_58536_54976# a_59097_54704# VSS sg13_lv_nmos ad=0.17p pd=1.68u as=0.17p ps=1.68u w=0.5u l=0.15u
X468 VSS a_56887_49467# VSS VSS sg13_lv_nmos ad=95f pd=0.88u as=0 ps=0 w=0.5u l=0.65u
X469 3bit_freq_divider_1.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 3bit_freq_divider_1.dff_nclk_0.nCLK VDD VDD sg13_lv_pmos ad=0.392p pd=2.94u as=0.392p ps=2.94u w=1.12u l=0.13u
X470 VSS a_52950_20401# 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.Q VSS sg13_lv_nmos ad=0.14505p pd=1.15u as=0.2516p ps=2.16u w=0.74u l=0.13u
X471 VSS vco_wob_0.vctl a_57112_40850# VSS sg13_lv_nmos ad=0.102p pd=1.28u as=65.99999f ps=0.74u w=0.3u l=0.13u
X472 a_62119_22361# a_61887_22290# a_61394_21976# VDD sg13_lv_pmos ad=79.8f pd=0.8u as=0.1428p ps=1.52u w=0.42u l=0.13u
X473 a_64383_23706# 3bit_freq_divider_1.dff_nclk_0.nRST VDD VDD sg13_lv_pmos ad=79.8f pd=0.8u as=79.8f ps=0.8u w=0.42u l=0.13u
X474 a_57111_40283# a_53022_43738# VDD VDD sg13_lv_pmos ad=59f pd=0.74u as=0.104p ps=1.34u w=0.2u l=0.13u
X475 a_51693_23426# a_51684_22692# a_51684_22284# VDD sg13_lv_pmos ad=79.8f pd=0.8u as=0.1428p ps=1.52u w=0.42u l=0.13u
X476 a_58454_40850# vco_wob_0.vctl VSS VSS sg13_lv_nmos ad=65.99999f pd=0.74u as=0.102p ps=1.28u w=0.3u l=0.13u
X477 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.nQ a_62654_20215# VDD VDD sg13_lv_pmos ad=0.7616p pd=3.6u as=0.2163p ps=1.55u w=1.12u l=0.13u
X478 VDD a_62654_21971# a_62900_21935# VDD sg13_lv_pmos ad=0.2163p pd=1.55u as=79.8f ps=0.8u w=0.42u l=0.13u
X479 a_54504_22015# 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.D a_55086_21975# VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=50.4f ps=0.66u w=0.42u l=0.13u
X480 a_55770_40850# a_55831_40413# a_54489_40413# VSS sg13_lv_nmos ad=0.17p pd=1.68u as=0.11p ps=0.94u w=0.5u l=0.13u
X481 a_54602_21487# 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.Q 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.D VSS sg13_lv_nmos ad=88.8f pd=0.98u as=0.1628p ps=1.18u w=0.74u l=0.13u
X482 a_56039_25022# a_56013_24979# a_55941_24882# VSS sg13_lv_nmos ad=0.2307p pd=1.615u as=0.27427p ps=2.28u w=0.795u l=0.13u
X483 a_51685_23725# a_51648_24041# a_52119_23843# VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=47.25f ps=0.645u w=0.42u l=0.13u
X484 a_54898_22885# 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.Q a_54434_23148# VDD sg13_lv_pmos ad=0.1225p pd=1.245u as=0.34p ps=2.68u w=1u l=0.13u
X485 a_51693_23426# a_51631_22774# a_51684_22284# VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0.1428p ps=1.52u w=0.42u l=0.13u
X486 VSS a_56887_49467# VSS VSS sg13_lv_nmos ad=95f pd=0.88u as=0 ps=0 w=0.5u l=0.65u
X487 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.D a_61707_21488# a_61878_21130# VDD sg13_lv_pmos ad=0.3808p pd=2.92u as=0.2128p ps=1.5u w=1.12u l=0.13u
X488 VSS 3bit_freq_divider_1.dff_nclk_0.sg13g2_dfrbp_1_0.CLK a_64383_23628# VSS sg13_lv_nmos ad=0.1544p pd=1.235u as=0.2516p ps=2.16u w=0.74u l=0.13u
X489 VSS 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.Q a_53054_24999# VSS sg13_lv_nmos ad=0.15245p pd=1.17u as=88.8f ps=0.98u w=0.74u l=0.13u
X490 a_61887_20534# a_61691_20534# VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0.19p ps=1.38u w=1u l=0.13u
X491 VSS a_56887_49467# VSS VSS sg13_lv_nmos ad=95f pd=0.88u as=0 ps=0 w=0.5u l=0.65u
X492 VSS a_56887_49467# VSS VSS sg13_lv_nmos ad=95f pd=0.88u as=0 ps=0 w=0.5u l=0.65u
X493 a_64714_21300# 3bit_freq_divider_1.sg13g2_or3_1_0.A VDD VDD sg13_lv_pmos ad=0.22p pd=1.44u as=0.3822p ps=1.84u w=1u l=0.13u
X494 a_54504_20259# 3bit_freq_divider_0.dff_nclk_0.nCLK VDD VDD sg13_lv_pmos ad=79.8f pd=0.8u as=0.1428p ps=1.52u w=0.42u l=0.13u
X495 a_61707_21488# 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.Q a_61675_21130# VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0.1225p ps=1.245u w=1u l=0.13u
X496 VDD 3bit_freq_divider_1.dff_nclk_0.sg13g2_dfrbp_1_0.CLK a_64383_23628# VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0.34p ps=2.68u w=1u l=0.13u
X497 a_51684_22692# a_51631_22774# VSS VSS sg13_lv_nmos ad=0.2516p pd=2.16u as=0.1544p ps=1.235u w=0.74u l=0.13u
X498 a_57111_40283# a_53022_43738# VDD VDD sg13_lv_pmos ad=59.75f pd=0.745u as=59f ps=0.74u w=0.2u l=0.13u
X499 a_57112_40850# a_57173_40413# a_55831_40413# VSS sg13_lv_nmos ad=0.17p pd=1.68u as=0.11p ps=0.94u w=0.5u l=0.13u
X500 VDD a_53774_20178# a_53738_20514# VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0.34p ps=2.68u w=1u l=0.13u
X501 VDD a_51693_23075# a_51729_23026# VDD sg13_lv_pmos ad=0.11785p pd=1.025u as=51.45f ps=0.665u w=0.42u l=0.13u
X502 VSS charge_pump_0.vout VSS VSS sg13_lv_nmos ad=0.285p pd=1.88u as=0 ps=0 w=1.5u l=0.65u
X503 a_45451_28860# CLK_IN a_45579_29803# VSS sg13_lv_nmos ad=68.39999f pd=0.74u as=68.39999f ps=0.74u w=0.36u l=0.15u
X504 a_55345_21385# 3bit_freq_divider_0.freq_div_cell_0.Cout a_55485_21477# VSS sg13_lv_nmos ad=0.2176p pd=1.96u as=0.1216p ps=1.02u w=0.64u l=0.13u
X505 a_57173_40413# a_58515_40413# a_58454_40850# VSS sg13_lv_nmos ad=0.11p pd=0.94u as=0.17p ps=1.68u w=0.5u l=0.13u
X506 charge_pump_0.bias_p charge_pump_0.bias_n a_56742_53480# VSS sg13_lv_nmos ad=0.34p pd=2.68u as=0.34p ps=2.68u w=1u l=1u
X507 VSS a_56887_49467# VSS VSS sg13_lv_nmos ad=95f pd=0.88u as=0 ps=0 w=0.5u l=0.65u
X508 a_62270_22299# a_62119_22361# VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0.34p ps=2.68u w=1u l=0.13u
X509 VSS a_56887_49467# VSS VSS sg13_lv_nmos ad=95f pd=0.88u as=0 ps=0 w=0.5u l=0.65u
X510 a_64817_23685# a_64383_23434# a_64383_23889# VDD sg13_lv_pmos ad=43.05f pd=0.625u as=0.17695p ps=1.56u w=0.42u l=0.13u
X511 a_51648_24041# a_51631_22774# a_51693_23075# VDD sg13_lv_pmos ad=0.17695p pd=1.56u as=0.19p ps=1.38u w=1u l=0.13u
X512 VDD a_45658_27900# PFD_0.DOWN VDD sg13_lv_pmos ad=60.8f pd=0.7u as=0.1088p ps=1.32u w=0.32u l=0.15u
X513 3bit_freq_divider_1.freq_div_cell_0.Cout a_60967_23234# VDD VDD sg13_lv_pmos ad=0.3808p pd=2.92u as=0.1918p ps=1.5u w=1.12u l=0.13u
X514 a_64419_23844# 3bit_freq_divider_1.dff_nclk_0.nRST VSS VSS sg13_lv_nmos ad=47.25f pd=0.645u as=90.3f ps=0.85u w=0.42u l=0.13u
X515 3bit_freq_divider_1.sg13g2_or3_1_0.C Y0 a_63520_25000# VSS sg13_lv_nmos ad=0.1628p pd=1.18u as=88.8f ps=0.98u w=0.74u l=0.13u
X516 VSS a_64383_23889# a_64384_24445# VSS sg13_lv_nmos ad=0.14505p pd=1.15u as=0.187p ps=1.78u w=0.55u l=0.13u
X517 a_64384_21091# 3bit_freq_divider_1.sg13g2_or3_1_0.C a_64714_21414# VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0.1275p ps=1.255u w=1u l=0.13u
X518 VSS charge_pump_0.vout VSS VSS sg13_lv_nmos ad=0.285p pd=1.88u as=0 ps=0 w=1.5u l=0.65u
X519 VSS a_53968_20434# a_53899_20488# VSS sg13_lv_nmos ad=0.1825p pd=1.325u as=0.19397p ps=1.29u w=0.64u l=0.13u
X520 a_45451_28860# CLK_IN a_45579_29803# VSS sg13_lv_nmos ad=68.39999f pd=0.74u as=68.39999f ps=0.74u w=0.36u l=0.15u
X521 VDD 3bit_freq_divider_1.dff_nclk_0.nCLK a_61394_20220# VDD sg13_lv_pmos ad=0.1428p pd=1.52u as=79.8f ps=0.8u w=0.42u l=0.13u
X522 a_54489_40413# VSS cap_cmim l=6.99u w=6.99u
X523 VSS a_53065_23691# 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.nQ VSS sg13_lv_nmos ad=0.2516p pd=2.16u as=0.2775p ps=2.23u w=0.74u l=0.13u
X524 a_53899_20488# a_53774_20178# a_53065_20179# VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0.17695p ps=1.56u w=1u l=0.13u
X525 a_52074_23129# a_51693_23075# a_52074_23051# VSS sg13_lv_nmos ad=48.3f pd=0.65u as=54.6f ps=0.68u w=0.42u l=0.13u
X526 a_62324_23772# a_62270_24055# a_62246_23772# VSS sg13_lv_nmos ad=48.3f pd=0.65u as=54.6f ps=0.68u w=0.42u l=0.13u
X527 VDD CLK_IN a_45579_29803# VDD sg13_lv_pmos ad=60.8f pd=0.7u as=0.1088p ps=1.32u w=0.32u l=0.15u
X528 a_54352_24116# a_53899_24000# VDD VDD sg13_lv_pmos ad=51.45f pd=0.665u as=0.11785p ps=1.025u w=0.42u l=0.13u
X529 VDD X1 a_52924_22885# VDD sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X530 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.D 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.Q a_61972_21488# VSS sg13_lv_nmos ad=0.1628p pd=1.18u as=88.8f ps=0.98u w=0.74u l=0.13u
X531 VDD 3bit_freq_divider_1.freq_div_cell_0.Cin a_61878_22886# VDD sg13_lv_pmos ad=0.2128p pd=1.5u as=0.3808p ps=2.92u w=1.12u l=0.13u
X532 VSS a_53774_23690# a_53738_24026# VSS sg13_lv_nmos ad=0.1544p pd=1.235u as=0.2516p ps=2.16u w=0.74u l=0.13u
X533 a_54489_40413# a_55831_40413# a_55769_40283# VDD sg13_lv_pmos ad=0.11p pd=0.94u as=0.17p ps=1.68u w=0.5u l=0.13u
X534 a_61061_23234# 3bit_freq_divider_1.freq_div_cell_0.Cin a_60967_23234# VSS sg13_lv_nmos ad=0.1216p pd=1.02u as=0.2176p ps=1.96u w=0.64u l=0.13u
X535 a_55862_56737# charge_pump_0.bias_p charge_pump_0.bias_n VDD sg13_lv_pmos ad=0.38p pd=2.38u as=0.68p ps=4.68u w=2u l=1u
X536 a_62900_21935# a_62654_21971# a_63038_21971# VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=47.25f ps=0.645u w=0.42u l=0.13u
X537 a_63038_21971# 3bit_freq_divider_1.dff_nclk_0.nCLK VSS VSS sg13_lv_nmos ad=47.25f pd=0.645u as=90.3f ps=0.85u w=0.42u l=0.13u
X538 VSS charge_pump_0.vout VSS VSS sg13_lv_nmos ad=0.285p pd=1.88u as=0 ps=0 w=1.5u l=0.65u
X539 3bit_freq_divider_0.dff_nclk_0.D a_51648_24041# VSS VSS sg13_lv_nmos ad=0.2775p pd=2.23u as=0.2516p ps=2.16u w=0.74u l=0.13u
X540 a_51721_24988# a_51721_24988# a_52065_24890# VSS sg13_lv_nmos ad=0.102p pd=1.28u as=0.2307p ps=1.615u w=0.3u l=0.13u
X541 VSS a_55345_23141# 3bit_freq_divider_0.freq_div_cell_0.Cout VSS sg13_lv_nmos ad=0.1331p pd=1.12u as=0.2516p ps=2.16u w=0.74u l=0.13u
X542 a_52886_24904# X0 VSS VSS sg13_lv_nmos ad=0.17462p pd=1.185u as=0.15245p ps=1.17u w=0.55u l=0.13u
X543 VSS charge_pump_0.vout VSS VSS sg13_lv_nmos ad=0.285p pd=1.88u as=0 ps=0 w=1.5u l=0.65u
X544 a_55831_40413# a_57173_40413# a_57111_40283# VDD sg13_lv_pmos ad=0.11p pd=0.94u as=0.17p ps=1.68u w=0.5u l=0.13u
X545 a_54504_23771# 3bit_freq_divider_0.dff_nclk_0.nCLK VDD VDD sg13_lv_pmos ad=79.8f pd=0.8u as=0.1428p ps=1.52u w=0.42u l=0.13u
X546 a_62119_24117# a_61691_24046# a_61394_23732# VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0.1428p ps=1.52u w=0.42u l=0.13u
X547 VSS 3bit_freq_divider_1.dff_nclk_0.nCLK a_61488_23732# VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=50.4f ps=0.66u w=0.42u l=0.13u
X548 3bit_freq_divider_0.EN nEN VSS VSS sg13_lv_nmos ad=0.259p pd=2.18u as=0.259p ps=2.18u w=0.74u l=0.13u
X549 VSS charge_pump_0.vout VSS VSS sg13_lv_nmos ad=0.285p pd=1.88u as=0 ps=0 w=1.5u l=0.65u
X550 a_59799_40285# a_53022_43738# VDD VDD sg13_lv_pmos ad=59.75f pd=0.745u as=59f ps=0.74u w=0.2u l=0.13u
X551 a_53899_20488# a_53738_20514# a_53065_20179# VSS sg13_lv_nmos ad=0.19397p pd=1.29u as=0.2017p ps=1.48u w=0.64u l=0.13u
X552 VSS PFD_0.VCO_CLK a_45451_28860# VSS sg13_lv_nmos ad=0.1224p pd=1.4u as=0.1224p ps=1.4u w=0.36u l=0.15u
X553 VSS a_46817_27899# a_45658_27900# VSS sg13_lv_nmos ad=0.1224p pd=1.4u as=0.1224p ps=1.4u w=0.36u l=0.15u
X554 a_53054_21487# X2 3bit_freq_divider_0.sg13g2_or3_1_0.A VSS sg13_lv_nmos ad=88.8f pd=0.98u as=0.1628p ps=1.18u w=0.74u l=0.13u
X555 a_53350_22885# X1 a_52886_23148# VDD sg13_lv_pmos ad=0.1225p pd=1.245u as=0.34p ps=2.68u w=1u l=0.13u
X556 VSS vco_wob_0.vctl a_57311_42591# VSS sg13_lv_nmos ad=0.102p pd=1.28u as=65.99999f ps=0.74u w=0.3u l=0.13u
X557 a_62900_23691# 3bit_freq_divider_1.dff_nclk_0.nCLK VDD VDD sg13_lv_pmos ad=79.8f pd=0.8u as=79.8f ps=0.8u w=0.42u l=0.13u
X558 a_53774_23690# 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.sg13g2_dfrbp_1_0.CLK VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0.19p ps=1.38u w=1u l=0.13u
X559 a_57311_42591# a_55836_43159# a_57178_43159# VSS sg13_lv_nmos ad=0.17p pd=1.68u as=0.11p ps=0.94u w=0.5u l=0.13u
X560 a_58653_42591# vco_wob_0.vctl VSS VSS sg13_lv_nmos ad=65.99999f pd=0.74u as=0.102p ps=1.28u w=0.3u l=0.13u
X561 a_55831_40413# a_57173_40413# a_57111_40283# VDD sg13_lv_pmos ad=0.1106p pd=0.945u as=0.11p ps=0.94u w=0.5u l=0.13u
X562 a_60967_21478# 3bit_freq_divider_1.freq_div_cell_0.Cout VDD VDD sg13_lv_pmos ad=0.1596p pd=1.22u as=0.2856p ps=2.36u w=0.84u l=0.13u
X563 VSS a_62900_21935# a_62848_21971# VSS sg13_lv_nmos ad=90.3f pd=0.85u as=54.6f ps=0.68u w=0.42u l=0.13u
X564 a_58426_43159# a_57178_43159# 3bit_freq_divider_0.CLK_IN VDD sg13_lv_pmos ad=0.17p pd=1.68u as=0.11p ps=0.94u w=0.5u l=0.13u
X565 3bit_freq_divider_0.CLK_IN a_57178_43159# a_58653_42591# VSS sg13_lv_nmos ad=0.11p pd=0.94u as=0.17p ps=1.68u w=0.5u l=0.13u
X566 VDD 3bit_freq_divider_0.dff_nclk_0.nCLK a_53968_20434# VDD sg13_lv_pmos ad=0.11785p pd=1.025u as=0.1533p ps=1.57u w=0.42u l=0.13u
X567 a_62119_24117# a_61887_24046# a_61394_23732# VDD sg13_lv_pmos ad=79.8f pd=0.8u as=0.1428p ps=1.52u w=0.42u l=0.13u
X568 a_54747_49259# charge_pump_0.bias_n VSS VSS sg13_lv_nmos ad=0.207p pd=1.545u as=0.408p ps=3.08u w=1.2u l=0.13u
X569 VDD a_53022_43738# a_54400_43159# VDD sg13_lv_pmos ad=59f pd=0.74u as=59.75f ps=0.745u w=0.2u l=0.13u
X570 VDD a_53022_43738# a_53022_43738# VDD sg13_lv_pmos ad=59f pd=0.74u as=59f ps=0.74u w=0.2u l=0.13u
X571 VSS 3bit_freq_divider_1.dff_nclk_0.nCLK a_62324_20260# VSS sg13_lv_nmos ad=0.1825p pd=1.325u as=48.3f ps=0.65u w=0.42u l=0.13u
X572 a_62848_21971# a_61691_22290# a_62654_21971# VSS sg13_lv_nmos ad=54.6f pd=0.68u as=0.2017p ps=1.48u w=0.42u l=0.13u
X573 a_63255_23244# Y1 a_63223_22886# VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0.1225p ps=1.245u w=1u l=0.13u
X574 a_53774_23690# 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.sg13g2_dfrbp_1_0.CLK VSS VSS sg13_lv_nmos ad=0.2516p pd=2.16u as=0.1544p ps=1.235u w=0.74u l=0.13u
X575 VSS 3bit_freq_divider_0.sg13g2_tiehi_1.L_HI a_54434_24904# VSS sg13_lv_nmos ad=0.374p pd=2.46u as=0.17462p ps=1.185u w=0.55u l=0.13u
X576 a_60385_24558# a_60385_24947# a_60385_24717# VDD sg13_lv_pmos ad=0.4657p pd=2.54u as=0.2442p ps=2.06u w=0.66u l=0.13u
X577 VSS Y1 a_63255_23244# VSS sg13_lv_nmos ad=0.15245p pd=1.17u as=0.17462p ps=1.185u w=0.55u l=0.13u
X578 a_58453_40283# a_58515_40413# a_57173_40413# VDD sg13_lv_pmos ad=0.17p pd=1.68u as=0.1106p ps=0.945u w=0.5u l=0.13u
X579 a_46749_30782# CLK_IN CLK_IN VDD sg13_lv_pmos ad=0.1088p pd=1.32u as=60.8f ps=0.7u w=0.32u l=0.15u
X580 a_61675_21130# 3bit_freq_divider_1.freq_div_cell_0.Cout VDD VDD sg13_lv_pmos ad=0.1225p pd=1.245u as=0.36p ps=2.72u w=1u l=0.13u
X581 a_52119_23653# a_51631_22774# a_51648_24041# VSS sg13_lv_nmos ad=54.6f pd=0.68u as=0.2017p ps=1.48u w=0.42u l=0.13u
X582 a_52950_22157# a_53065_21935# VDD VDD sg13_lv_pmos ad=0.2856p pd=2.36u as=0.2016p ps=1.5u w=0.84u l=0.13u
X583 PFD_0.VCO_CLK a_51648_24438# VDD VDD sg13_lv_pmos ad=0.3808p pd=2.92u as=0.2016p ps=1.5u w=1.12u l=0.13u
X584 3bit_freq_divider_1.dff_nclk_0.D a_64383_23889# VSS VSS sg13_lv_nmos ad=0.2775p pd=2.23u as=0.2516p ps=2.16u w=0.74u l=0.13u
X585 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 3bit_freq_divider_1.sg13g2_nand2_1_0.Y VDD VDD sg13_lv_pmos ad=0.392p pd=2.94u as=0.392p ps=2.94u w=1.12u l=0.13u
X586 VDD a_62900_20179# a_62879_20613# VDD sg13_lv_pmos ad=79.8f pd=0.8u as=43.05f ps=0.625u w=0.42u l=0.13u
X587 a_55345_21385# 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.Q VDD VDD sg13_lv_pmos ad=0.1596p pd=1.22u as=0.1918p ps=1.5u w=0.84u l=0.13u
X588 VDD a_53065_20179# 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.nQ VDD sg13_lv_pmos ad=0.2163p pd=1.55u as=0.7616p ps=3.6u w=1.12u l=0.13u
X589 a_51648_21103# 3bit_freq_divider_0.sg13g2_or3_1_0.A VSS VSS sg13_lv_nmos ad=0.198p pd=1.27u as=0.13395p ps=1.12u w=0.55u l=0.13u
X590 VSS a_51648_21103# 3bit_freq_divider_0.dff_nclk_0.nCLK VSS sg13_lv_nmos ad=0.13395p pd=1.12u as=0.2516p ps=2.16u w=0.74u l=0.13u
X591 a_52944_43077# a_53147_40413# a_53085_40283# VDD sg13_lv_pmos ad=0.1106p pd=0.945u as=0.11p ps=0.94u w=0.5u l=0.13u
X592 a_59799_40285# 3bit_freq_divider_0.CLK_IN a_58515_40413# VDD sg13_lv_pmos ad=0.11p pd=0.94u as=0.11p ps=0.94u w=0.5u l=0.13u
X593 a_53065_23691# a_53738_24026# a_53702_24124# VDD sg13_lv_pmos ad=0.17695p pd=1.56u as=43.05f ps=0.625u w=0.42u l=0.13u
X594 a_54504_22015# a_53738_22270# a_53968_22190# VDD sg13_lv_pmos ad=0.1428p pd=1.52u as=79.8f ps=0.8u w=0.42u l=0.13u
X595 VDD a_53022_43738# a_54400_43159# VDD sg13_lv_pmos ad=0.104p pd=1.34u as=59f ps=0.74u w=0.2u l=0.13u
X596 VDD a_62654_21971# a_63463_21972# VDD sg13_lv_pmos ad=0.2016p pd=1.5u as=0.2856p ps=2.36u w=0.84u l=0.13u
X597 a_47954_28913# PFD_0.VCO_CLK VDD VDD sg13_lv_pmos ad=0.1088p pd=1.32u as=60.8f ps=0.7u w=0.32u l=0.15u
X598 VDD 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.Q a_60967_24990# VDD sg13_lv_pmos ad=0.1918p pd=1.5u as=0.1596p ps=1.22u w=0.84u l=0.13u
X599 a_52950_20401# a_53065_20179# VSS VSS sg13_lv_nmos ad=0.187p pd=1.78u as=0.14505p ps=1.15u w=0.55u l=0.13u
X600 a_53086_40850# vco_wob_0.vctl VSS VSS sg13_lv_nmos ad=65.99999f pd=0.74u as=0.102p ps=1.28u w=0.3u l=0.13u
X601 a_62246_23772# a_61887_24046# a_62119_24117# VSS sg13_lv_nmos ad=54.6f pd=0.68u as=79.8f ps=0.8u w=0.42u l=0.13u
X602 VDD 3bit_freq_divider_0.freq_div_cell_0.Cin a_54898_22885# VDD sg13_lv_pmos ad=0.36p pd=2.72u as=0.1225p ps=1.245u w=1u l=0.13u
X603 VDD a_53022_43738# a_57111_40283# VDD sg13_lv_pmos ad=0.104p pd=1.34u as=59.75f ps=0.745u w=0.2u l=0.13u
X604 a_48909_28913# PFD_0.VCO_CLK a_47954_28913# VSS sg13_lv_nmos ad=68.39999f pd=0.74u as=68.39999f ps=0.74u w=0.36u l=0.15u
X605 VSS 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.Q a_52886_21392# VSS sg13_lv_nmos ad=0.374p pd=2.46u as=0.17462p ps=1.185u w=0.55u l=0.13u
X606 a_55345_24897# 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.Q VDD VDD sg13_lv_pmos ad=0.1596p pd=1.22u as=0.1918p ps=1.5u w=0.84u l=0.13u
X607 VSS charge_pump_0.vout VSS VSS sg13_lv_nmos ad=0.285p pd=1.88u as=0 ps=0 w=1.5u l=0.65u
X608 a_58453_40283# a_53022_43738# VDD VDD sg13_lv_pmos ad=59.75f pd=0.745u as=59f ps=0.74u w=0.2u l=0.13u
X609 3bit_freq_divider_0.sg13g2_or3_1_0.B a_52886_23148# VSS VSS sg13_lv_nmos ad=0.1628p pd=1.18u as=0.3108p ps=2.32u w=0.74u l=0.13u
X610 VSS a_62654_20215# a_63463_20216# VSS sg13_lv_nmos ad=0.14505p pd=1.15u as=0.187p ps=1.78u w=0.55u l=0.13u
X611 a_63255_21488# 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.Q VSS VSS sg13_lv_nmos ad=0.17462p pd=1.185u as=0.374p ps=2.46u w=0.55u l=0.13u
X612 a_54252_22015# 3bit_freq_divider_0.dff_nclk_0.nCLK VSS VSS sg13_lv_nmos ad=48.3f pd=0.65u as=0.1825p ps=1.325u w=0.42u l=0.13u
X613 a_63426_22886# Y1 VDD VDD sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X614 VDD a_53022_43738# a_55742_43159# VDD sg13_lv_pmos ad=0.104p pd=1.34u as=59f ps=0.74u w=0.2u l=0.13u
X615 a_51685_23725# 3bit_freq_divider_0.dff_nclk_0.nRST VDD VDD sg13_lv_pmos ad=79.8f pd=0.8u as=79.8f ps=0.8u w=0.42u l=0.13u
X616 a_53539_20214# a_53065_20179# a_53445_20214# VSS sg13_lv_nmos ad=47.25f pd=0.645u as=0.1428p ps=1.52u w=0.42u l=0.13u
X617 VSS 3bit_freq_divider_0.dff_nclk_0.nCLK a_53539_20214# VSS sg13_lv_nmos ad=90.3f pd=0.85u as=47.25f ps=0.645u w=0.42u l=0.13u
X618 VDD 3bit_freq_divider_0.EN 3bit_freq_divider_0.sg13g2_nand2_1_0.Y VDD sg13_lv_pmos ad=0.3808p pd=2.92u as=0.2128p ps=1.5u w=1.12u l=0.13u
X619 a_54504_22015# a_53774_21934# a_53968_22190# VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=79.8f ps=0.8u w=0.42u l=0.13u
X620 3bit_freq_divider_1.sg13g2_or3_1_0.A a_63255_21488# a_63426_21130# VDD sg13_lv_pmos ad=0.3808p pd=2.92u as=0.2128p ps=1.5u w=1.12u l=0.13u
X621 a_52924_21129# a_52886_21392# 3bit_freq_divider_0.sg13g2_or3_1_0.A VDD sg13_lv_pmos ad=0.2128p pd=1.5u as=0.3808p ps=2.92u w=1.12u l=0.13u
X622 VDD 3bit_freq_divider_1.dff_nclk_0.nCLK a_61394_21976# VDD sg13_lv_pmos ad=0.1428p pd=1.52u as=79.8f ps=0.8u w=0.42u l=0.13u
X623 a_57178_43159# a_55836_43159# a_57084_43159# VDD sg13_lv_pmos ad=0.11p pd=0.94u as=0.11p ps=0.94u w=0.5u l=0.13u
X624 VSS 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.sg13g2_dfrbp_1_0.CLK a_61691_20534# VSS sg13_lv_nmos ad=0.1544p pd=1.235u as=0.2516p ps=2.16u w=0.74u l=0.13u
X625 a_53968_20434# a_53774_20178# a_54352_20604# VDD sg13_lv_pmos ad=79.8f pd=0.8u as=51.45f ps=0.665u w=0.42u l=0.13u
X626 a_64419_23326# a_64383_23300# VSS VSS sg13_lv_nmos ad=0.19397p pd=1.29u as=0.1825p ps=1.325u w=0.64u l=0.13u
X627 a_52944_43077# a_53147_40413# a_53086_40850# VSS sg13_lv_nmos ad=0.11p pd=0.94u as=0.17p ps=1.68u w=0.5u l=0.13u
X628 3bit_freq_divider_1.sg13g2_nand2_1_0.Y 3bit_freq_divider_0.EN VDD VDD sg13_lv_pmos ad=0.2128p pd=1.5u as=0.3808p ps=2.92u w=1.12u l=0.13u
X629 VSS charge_pump_0.vout VSS VSS sg13_lv_nmos ad=0.285p pd=1.88u as=0 ps=0 w=1.5u l=0.65u
X630 a_47954_28913# PFD_0.VCO_CLK a_46817_27899# VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0.1428p ps=1.52u w=0.42u l=0.15u
X631 a_62270_22299# a_62119_22361# VSS VSS sg13_lv_nmos ad=0.19397p pd=1.29u as=0.1825p ps=1.325u w=0.64u l=0.13u
X632 a_62900_23691# a_62654_23727# a_63038_23727# VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=47.25f ps=0.645u w=0.42u l=0.13u
X633 a_63038_23727# 3bit_freq_divider_1.dff_nclk_0.nCLK VSS VSS sg13_lv_nmos ad=47.25f pd=0.645u as=90.3f ps=0.85u w=0.42u l=0.13u
X634 VDD a_53022_43738# a_53022_43738# VDD sg13_lv_pmos ad=0.104p pd=1.34u as=59.75f ps=0.745u w=0.2u l=0.13u
X635 a_52924_24641# a_52886_24904# 3bit_freq_divider_0.sg13g2_or3_1_0.C VDD sg13_lv_pmos ad=0.2128p pd=1.5u as=0.3808p ps=2.92u w=1.12u l=0.13u
X636 a_56137_24678# a_56137_24678# a_56039_25022# VSS sg13_lv_nmos ad=0.102p pd=1.28u as=0.2307p ps=1.615u w=0.3u l=0.13u
X637 a_45579_29803# CLK_IN a_45451_28860# VSS sg13_lv_nmos ad=68.39999f pd=0.74u as=0.1224p ps=1.4u w=0.36u l=0.15u
X638 VSS a_45658_27900# PFD_0.DOWN VSS sg13_lv_nmos ad=0.1632p pd=1.64u as=0.1632p ps=1.64u w=0.48u l=0.15u
X639 a_52944_43077# VSS cap_cmim l=6.99u w=6.99u
X640 a_53702_22368# a_53445_21970# VDD VDD sg13_lv_pmos ad=43.05f pd=0.625u as=79.8f ps=0.8u w=0.42u l=0.13u
X641 a_63520_23244# 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.Q VSS VSS sg13_lv_nmos ad=88.8f pd=0.98u as=0.15245p ps=1.17u w=0.74u l=0.13u
X642 a_61707_23244# 3bit_freq_divider_1.freq_div_cell_0.Cin VSS VSS sg13_lv_nmos ad=0.17462p pd=1.185u as=0.374p ps=2.46u w=0.55u l=0.13u
X643 a_51759_25014# a_51721_24988# a_51600_24907# VDD sg13_lv_pmos ad=0.2442p pd=2.06u as=0.4657p ps=2.54u w=0.66u l=0.13u
X644 VDD a_53968_23946# a_53899_24000# VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0.19p ps=1.38u w=1u l=0.13u
X645 VDD 3bit_freq_divider_0.freq_div_cell_0.Cout a_55345_21385# VDD sg13_lv_pmos ad=0.2856p pd=2.36u as=0.1596p ps=1.22u w=0.84u l=0.13u
X646 VSS 3bit_freq_divider_0.freq_div_cell_0.Cout a_54602_21487# VSS sg13_lv_nmos ad=0.15245p pd=1.17u as=88.8f ps=0.98u w=0.74u l=0.13u
X647 VSS a_56887_49467# VSS VSS sg13_lv_nmos ad=95f pd=0.88u as=0 ps=0 w=0.5u l=0.65u
X648 a_53058_43159# a_53022_43738# VDD VDD sg13_lv_pmos ad=59f pd=0.74u as=59f ps=0.74u w=0.2u l=0.13u
X649 VSS a_64384_21091# 3bit_freq_divider_1.dff_nclk_0.nCLK VSS sg13_lv_nmos ad=0.13395p pd=1.12u as=0.2516p ps=2.16u w=0.74u l=0.13u
X650 VDD a_62270_22299# a_62221_22361# VDD sg13_lv_pmos ad=0.11785p pd=1.025u as=51.45f ps=0.665u w=0.42u l=0.13u
X651 VSS vco_wob_0.vctl a_54627_42591# VSS sg13_lv_nmos ad=0.102p pd=1.28u as=65.99999f ps=0.74u w=0.3u l=0.13u
X652 a_51721_23684# a_51684_22692# a_51648_24041# VDD sg13_lv_pmos ad=43.05f pd=0.625u as=0.17695p ps=1.56u w=0.42u l=0.13u
X653 a_54627_42591# a_53152_43159# a_54494_43159# VSS sg13_lv_nmos ad=0.17p pd=1.68u as=0.11p ps=0.94u w=0.5u l=0.13u
X654 a_51684_22284# 3bit_freq_divider_0.dff_nclk_0.D VDD VDD sg13_lv_pmos ad=79.8f pd=0.8u as=0.1428p ps=1.52u w=0.42u l=0.13u
X655 a_61887_24046# a_61691_24046# VSS VSS sg13_lv_nmos ad=0.2516p pd=2.16u as=0.1544p ps=1.235u w=0.74u l=0.13u
X656 VDD a_53065_23691# 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.nQ VDD sg13_lv_pmos ad=0.2163p pd=1.55u as=0.7616p ps=3.6u w=1.12u l=0.13u
X657 a_53445_20214# a_53065_20179# VDD VDD sg13_lv_pmos ad=79.8f pd=0.8u as=0.2163p ps=1.55u w=0.42u l=0.13u
X658 VSS a_56887_49467# VSS VSS sg13_lv_nmos ad=95f pd=0.88u as=0 ps=0 w=0.5u l=0.65u
X659 VDD 3bit_freq_divider_0.sg13g2_tiehi_1.L_HI a_55345_24897# VDD sg13_lv_pmos ad=0.2856p pd=2.36u as=0.1596p ps=1.22u w=0.84u l=0.13u
X660 3bit_freq_divider_1.sg13g2_or3_1_0.A Y2 a_63520_21488# VSS sg13_lv_nmos ad=0.1628p pd=1.18u as=88.8f ps=0.98u w=0.74u l=0.13u
X661 VDD 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.Q a_54472_22885# VDD sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X662 CLK_OUT a_64384_24445# VDD VDD sg13_lv_pmos ad=0.3808p pd=2.92u as=0.2016p ps=1.5u w=1.12u l=0.13u
X663 VSS a_56887_49467# VSS VSS sg13_lv_nmos ad=95f pd=0.88u as=0 ps=0 w=0.5u l=0.65u
X664 a_53065_20179# a_53774_20178# a_53722_20214# VSS sg13_lv_nmos ad=0.2017p pd=1.48u as=54.6f ps=0.68u w=0.42u l=0.13u
X665 a_64424_22200# 3bit_freq_divider_1.dff_nclk_0.D VDD VDD sg13_lv_pmos ad=79.8f pd=0.8u as=0.1428p ps=1.52u w=0.42u l=0.13u
X666 a_63223_22886# 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.Q VDD VDD sg13_lv_pmos ad=0.1225p pd=1.245u as=0.36p ps=2.72u w=1u l=0.13u
X667 a_61488_21976# 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.D a_61394_21976# VSS sg13_lv_nmos ad=50.4f pd=0.66u as=0.1428p ps=1.52u w=0.42u l=0.13u
X668 VSS a_62900_23691# a_62848_23727# VSS sg13_lv_nmos ad=90.3f pd=0.85u as=54.6f ps=0.68u w=0.42u l=0.13u
X669 a_53722_20214# a_53445_20214# VSS VSS sg13_lv_nmos ad=54.6f pd=0.68u as=90.3f ps=0.85u w=0.42u l=0.13u
X670 a_64383_23706# a_64383_23889# a_64419_23844# VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=47.25f ps=0.645u w=0.42u l=0.13u
X671 VSS 3bit_freq_divider_1.dff_nclk_0.nCLK a_62324_22016# VSS sg13_lv_nmos ad=0.1825p pd=1.325u as=48.3f ps=0.65u w=0.42u l=0.13u
X672 a_62848_23727# a_61691_24046# a_62654_23727# VSS sg13_lv_nmos ad=54.6f pd=0.68u as=0.2017p ps=1.48u w=0.42u l=0.13u
X673 VDD charge_pump_0.bias_p a_54842_49733# VDD sg13_lv_pmos ad=0.1005p pd=1.34u as=55.5f ps=0.74u w=0.15u l=0.13u
X674 VSS a_56887_49467# VSS VSS sg13_lv_nmos ad=95f pd=0.88u as=0 ps=0 w=0.5u l=0.65u
X675 a_46817_27899# PFD_0.VCO_CLK PFD_0.VCO_CLK VDD sg13_lv_pmos ad=0.1088p pd=1.32u as=60.8f ps=0.7u w=0.32u l=0.15u
X676 a_57173_40413# a_58515_40413# a_58453_40283# VDD sg13_lv_pmos ad=0.1106p pd=0.945u as=0.11p ps=0.94u w=0.5u l=0.13u
X677 a_64384_21091# 3bit_freq_divider_1.sg13g2_or3_1_0.C VSS VSS sg13_lv_nmos ad=0.187p pd=1.78u as=0.1045p ps=0.93u w=0.55u l=0.13u
X678 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 3bit_freq_divider_1.sg13g2_nand2_1_0.Y VSS VSS sg13_lv_nmos ad=0.259p pd=2.18u as=0.259p ps=2.18u w=0.74u l=0.13u
X679 VSS charge_pump_0.vout VSS VSS sg13_lv_nmos ad=0.51p pd=3.68u as=0 ps=0 w=1.5u l=0.65u
X680 a_53285_42591# vco_wob_0.vctl VSS VSS sg13_lv_nmos ad=65.99999f pd=0.74u as=0.102p ps=1.28u w=0.3u l=0.13u
X681 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.D a_54434_24904# VSS VSS sg13_lv_nmos ad=0.1628p pd=1.18u as=0.3108p ps=2.32u w=0.74u l=0.13u
X682 a_54504_23771# a_53738_24026# a_53968_23946# VDD sg13_lv_pmos ad=0.1428p pd=1.52u as=79.8f ps=0.8u w=0.42u l=0.13u
X683 a_61878_22886# 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.Q VDD VDD sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X684 CLK_IN CLK_IN a_46749_30782# VDD sg13_lv_pmos ad=60.8f pd=0.7u as=0.1088p ps=1.32u w=0.32u l=0.15u
X685 a_53058_43159# a_52944_43077# a_53152_43159# VDD sg13_lv_pmos ad=0.17p pd=1.68u as=0.11p ps=0.94u w=0.5u l=0.13u
X686 a_53152_43159# a_52944_43077# a_53285_42591# VSS sg13_lv_nmos ad=0.11p pd=0.94u as=0.17p ps=1.68u w=0.5u l=0.13u
X687 a_54434_21392# 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.Q VSS VSS sg13_lv_nmos ad=0.17462p pd=1.185u as=0.15245p ps=1.17u w=0.55u l=0.13u
X688 VSS a_63255_25000# 3bit_freq_divider_1.sg13g2_or3_1_0.C VSS sg13_lv_nmos ad=0.3108p pd=2.32u as=0.1628p ps=1.18u w=0.74u l=0.13u
X689 a_47954_28913# PFD_0.VCO_CLK a_48909_28913# VSS sg13_lv_nmos ad=68.39999f pd=0.74u as=68.39999f ps=0.74u w=0.36u l=0.15u
X690 VDD 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.Q a_63426_24642# VDD sg13_lv_pmos ad=0.2128p pd=1.5u as=0.3808p ps=2.92u w=1.12u l=0.13u
X691 3bit_freq_divider_1.freq_div_cell_1.Cout a_60967_21478# VSS VSS sg13_lv_nmos ad=0.2516p pd=2.16u as=0.1331p ps=1.12u w=0.74u l=0.13u
X692 a_53085_40283# a_53147_40413# a_52944_43077# VDD sg13_lv_pmos ad=0.17p pd=1.68u as=0.1106p ps=0.945u w=0.5u l=0.13u
X693 a_54472_22885# 3bit_freq_divider_0.freq_div_cell_0.Cin VDD VDD sg13_lv_pmos ad=0.3808p pd=2.92u as=0.2128p ps=1.5u w=1.12u l=0.13u
X694 VSS charge_pump_0.vout VSS VSS sg13_lv_nmos ad=0.285p pd=1.88u as=0 ps=0 w=1.5u l=0.65u
X695 a_64383_23300# 3bit_freq_divider_1.dff_nclk_0.nRST VDD VDD sg13_lv_pmos ad=0.1533p pd=1.57u as=0.11785p ps=1.025u w=0.42u l=0.13u
X696 a_55769_40283# a_55831_40413# a_54489_40413# VDD sg13_lv_pmos ad=0.11p pd=0.94u as=0.11p ps=0.94u w=0.5u l=0.13u
X697 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.Q a_63463_21972# VSS VSS sg13_lv_nmos ad=0.2516p pd=2.16u as=0.14505p ps=1.15u w=0.74u l=0.13u
X698 a_54428_40850# vco_wob_0.vctl VSS VSS sg13_lv_nmos ad=65.99999f pd=0.74u as=0.102p ps=1.28u w=0.3u l=0.13u
X699 VDD PFD_0.VCO_CLK a_47954_28913# VDD sg13_lv_pmos ad=60.8f pd=0.7u as=0.1088p ps=1.32u w=0.32u l=0.15u
X700 a_54352_20604# a_53899_20488# VDD VDD sg13_lv_pmos ad=51.45f pd=0.665u as=0.11785p ps=1.025u w=0.42u l=0.13u
X701 charge_pump_0.vout a_56887_49467# rhigh l=0.96u w=0.5u
X702 a_55836_43159# a_54494_43159# a_55742_43159# VDD sg13_lv_pmos ad=0.11p pd=0.94u as=0.11p ps=0.94u w=0.5u l=0.13u
X703 VDD a_53022_43738# a_58453_40283# VDD sg13_lv_pmos ad=0.104p pd=1.34u as=59.75f ps=0.745u w=0.2u l=0.13u
X704 3bit_freq_divider_1.freq_div_cell_0.Cin a_60967_24990# VSS VSS sg13_lv_nmos ad=0.2516p pd=2.16u as=0.1331p ps=1.12u w=0.74u l=0.13u
X705 VSS 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.Q a_53054_21487# VSS sg13_lv_nmos ad=0.15245p pd=1.17u as=88.8f ps=0.98u w=0.74u l=0.13u
X706 VSS 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK a_61691_22290# VSS sg13_lv_nmos ad=0.1544p pd=1.235u as=0.2516p ps=2.16u w=0.74u l=0.13u
X707 VDD 3bit_freq_divider_0.dff_nclk_0.nCLK a_53445_23726# VDD sg13_lv_pmos ad=79.8f pd=0.8u as=79.8f ps=0.8u w=0.42u l=0.13u
X708 VSS charge_pump_0.vout VSS VSS sg13_lv_nmos ad=0.285p pd=1.88u as=0 ps=0 w=1.5u l=0.65u
X709 a_54472_21129# a_54434_21392# 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.D VDD sg13_lv_pmos ad=0.2128p pd=1.5u as=0.3808p ps=2.92u w=1.12u l=0.13u
X710 VDD 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.Q a_53350_21129# VDD sg13_lv_pmos ad=0.36p pd=2.72u as=0.1225p ps=1.245u w=1u l=0.13u
X711 a_57111_40283# a_57173_40413# a_55831_40413# VDD sg13_lv_pmos ad=0.11p pd=0.94u as=0.11p ps=0.94u w=0.5u l=0.13u
X712 a_52065_24890# a_51759_25014# a_51622_24863# VSS sg13_lv_nmos ad=0.2307p pd=1.615u as=0.27427p ps=2.28u w=0.795u l=0.13u
X713 a_62270_24055# a_62119_24117# VSS VSS sg13_lv_nmos ad=0.19397p pd=1.29u as=0.1825p ps=1.325u w=0.64u l=0.13u
X714 a_58426_43159# a_53022_43738# VDD VDD sg13_lv_pmos ad=59f pd=0.74u as=59f ps=0.74u w=0.2u l=0.13u
X715 a_57173_40413# a_58515_40413# a_58453_40283# VDD sg13_lv_pmos ad=0.11p pd=0.94u as=0.17p ps=1.68u w=0.5u l=0.13u
X716 VDD a_53022_43738# a_59799_40285# VDD sg13_lv_pmos ad=59f pd=0.74u as=59f ps=0.74u w=0.2u l=0.13u
X717 a_64383_23889# a_64383_23434# a_64419_23326# VSS sg13_lv_nmos ad=0.2017p pd=1.48u as=0.19397p ps=1.29u w=0.64u l=0.13u
X718 a_53085_40283# a_53022_43738# VDD VDD sg13_lv_pmos ad=59.75f pd=0.745u as=59f ps=0.74u w=0.2u l=0.13u
X719 VDD a_53022_43738# a_54427_40283# VDD sg13_lv_pmos ad=59f pd=0.74u as=59f ps=0.74u w=0.2u l=0.13u
X720 VDD a_53022_43738# a_59799_40285# VDD sg13_lv_pmos ad=0.104p pd=1.34u as=59.75f ps=0.745u w=0.2u l=0.13u
X721 a_62221_22361# a_61691_22290# a_62119_22361# VDD sg13_lv_pmos ad=51.45f pd=0.665u as=79.8f ps=0.8u w=0.42u l=0.13u
X722 a_56742_53480# VSS rhigh l=12u w=1u
X723 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.Q a_63463_23728# VDD VDD sg13_lv_pmos ad=0.3808p pd=2.92u as=0.2016p ps=1.5u w=1.12u l=0.13u
X724 a_53147_40413# a_54489_40413# a_54428_40850# VSS sg13_lv_nmos ad=0.11p pd=0.94u as=0.17p ps=1.68u w=0.5u l=0.13u
X725 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.D a_61707_23244# a_61878_22886# VDD sg13_lv_pmos ad=0.3808p pd=2.92u as=0.2128p ps=1.5u w=1.12u l=0.13u
X726 VDD a_62270_24055# a_62221_24117# VDD sg13_lv_pmos ad=0.11785p pd=1.025u as=51.45f ps=0.665u w=0.42u l=0.13u
X727 VSS charge_pump_0.vout VSS VSS sg13_lv_nmos ad=0.285p pd=1.88u as=0 ps=0 w=1.5u l=0.65u
X728 a_54472_24641# a_54434_24904# 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.D VDD sg13_lv_pmos ad=0.2128p pd=1.5u as=0.3808p ps=2.92u w=1.12u l=0.13u
X729 VDD 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.Q a_53350_24641# VDD sg13_lv_pmos ad=0.36p pd=2.72u as=0.1225p ps=1.245u w=1u l=0.13u
X730 a_53058_43159# a_52944_43077# a_53152_43159# VDD sg13_lv_pmos ad=0.11p pd=0.94u as=0.1106p ps=0.945u w=0.5u l=0.13u
X731 VDD 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.D a_54504_20259# VDD sg13_lv_pmos ad=0.1428p pd=1.52u as=79.8f ps=0.8u w=0.42u l=0.13u
X732 a_61707_23244# 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.Q a_61675_22886# VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0.1225p ps=1.245u w=1u l=0.13u
X733 a_64419_23326# a_64383_23300# VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0.34p ps=2.68u w=1u l=0.13u
X734 a_51708_21413# 3bit_freq_divider_0.sg13g2_or3_1_0.B a_51708_21299# VDD sg13_lv_pmos ad=0.1275p pd=1.255u as=0.22p ps=1.44u w=1u l=0.13u
X735 VSS 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.Q a_61707_23244# VSS sg13_lv_nmos ad=0.15245p pd=1.17u as=0.17462p ps=1.185u w=0.55u l=0.13u
X736 VSS a_53065_20179# 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.nQ VSS sg13_lv_nmos ad=0.2516p pd=2.16u as=0.2775p ps=2.23u w=0.74u l=0.13u
X737 a_62324_20260# a_62270_20543# a_62246_20260# VSS sg13_lv_nmos ad=48.3f pd=0.65u as=54.6f ps=0.68u w=0.42u l=0.13u
X738 a_62900_20179# 3bit_freq_divider_1.dff_nclk_0.nCLK VDD VDD sg13_lv_pmos ad=79.8f pd=0.8u as=79.8f ps=0.8u w=0.42u l=0.13u
X739 a_55836_43159# VSS cap_cmim l=6.99u w=6.99u
X740 a_53774_20178# 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.sg13g2_dfrbp_1_0.CLK VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0.19p ps=1.38u w=1u l=0.13u
X741 VSS a_53774_20178# a_53738_20514# VSS sg13_lv_nmos ad=0.1544p pd=1.235u as=0.2516p ps=2.16u w=0.74u l=0.13u
X742 VDD a_53022_43738# a_55742_43159# VDD sg13_lv_pmos ad=59f pd=0.74u as=59.75f ps=0.745u w=0.2u l=0.13u
X743 a_45579_29803# CLK_IN a_46749_30782# VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0.1428p ps=1.52u w=0.42u l=0.15u
X744 a_62119_20605# a_61887_20534# a_61394_20220# VDD sg13_lv_pmos ad=79.8f pd=0.8u as=0.1428p ps=1.52u w=0.42u l=0.13u
X745 a_62654_21971# a_61691_22290# a_62270_22299# VDD sg13_lv_pmos ad=0.17695p pd=1.56u as=0.19p ps=1.38u w=1u l=0.13u
X746 a_60479_25023# a_60385_24947# a_60385_24947# VSS sg13_lv_nmos ad=0.2307p pd=1.615u as=0.102p ps=1.28u w=0.3u l=0.13u
X747 a_64809_23027# a_64383_23628# a_64383_23300# VDD sg13_lv_pmos ad=51.45f pd=0.665u as=79.8f ps=0.8u w=0.42u l=0.13u
X748 3bit_freq_divider_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 3bit_freq_divider_0.dff_nclk_0.nCLK VSS VSS sg13_lv_nmos ad=0.259p pd=2.18u as=0.259p ps=2.18u w=0.74u l=0.13u
X749 a_64419_23654# a_64383_23628# a_64383_23889# VSS sg13_lv_nmos ad=54.6f pd=0.68u as=0.2017p ps=1.48u w=0.42u l=0.13u
X750 VSS vco_wob_0.vctl VSS VSS sg13_lv_nmos ad=0.1005p pd=1.34u as=0 ps=0 w=0.15u l=0.13u
X751 a_52886_21392# X2 VSS VSS sg13_lv_nmos ad=0.17462p pd=1.185u as=0.15245p ps=1.17u w=0.55u l=0.13u
X752 a_58536_54976# charge_pump_0.bias_n VSS VSS sg13_lv_nmos ad=0.34p pd=2.68u as=0.34p ps=2.68u w=1u l=1u
X753 VSS a_61707_25000# 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.D VSS sg13_lv_nmos ad=0.3108p pd=2.32u as=0.1628p ps=1.18u w=0.74u l=0.13u
X754 VDD a_53022_43738# a_57084_43159# VDD sg13_lv_pmos ad=59f pd=0.74u as=59.75f ps=0.745u w=0.2u l=0.13u
X755 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.nQ a_62654_21971# VDD VDD sg13_lv_pmos ad=0.7616p pd=3.6u as=0.2163p ps=1.55u w=1.12u l=0.13u
X756 VDD 3bit_freq_divider_0.sg13g2_nand2_1_0.Y 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.sg13g2_dfrbp_1_0.CLK VDD sg13_lv_pmos ad=0.392p pd=2.94u as=0.392p ps=2.94u w=1.12u l=0.13u
X757 VSS charge_pump_0.vout VSS VSS sg13_lv_nmos ad=0.285p pd=1.88u as=0 ps=0 w=1.5u l=0.65u
C0 a_60385_24717# VDD 0.11381f
C1 3bit_freq_divider_1.dff_nclk_0.nRST a_64383_23706# 0.25925f
C2 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.Q 3bit_freq_divider_0.sg13g2_or3_1_0.C 0.05745f
C3 3bit_freq_divider_1.dff_nclk_0.nCLK 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.D 0.21745f
C4 3bit_freq_divider_0.freq_div_cell_0.Cin a_55345_23141# 0.13034f
C5 a_64383_23706# a_64383_23434# 0.04306f
C6 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.Q a_63255_21488# 0.12248f
C7 3bit_freq_divider_1.dff_nclk_0.nCLK a_61691_22290# 0.35569f
C8 3bit_freq_divider_1.dff_nclk_0.nCLK a_62270_24055# 0.17312f
C9 a_53738_20514# a_53899_20488# 0.66077f
C10 charge_pump_0.bias_n VDD 0.83592f
C11 3bit_freq_divider_0.dff_nclk_0.nCLK a_53738_22270# 0.18642f
C12 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.Q Y2 0.21293f
C13 a_53065_21935# 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.Q 0.0119f
C14 charge_pump_0.bias_n PFD_0.DOWN 0.01578f
C15 a_54489_40413# VDD 1.15543f
C16 a_51684_22284# VDD 0.36995f
C17 3bit_freq_divider_1.freq_div_cell_0.Cin 3bit_freq_divider_1.sg13g2_nand2_1_0.Y 0.25573f
C18 3bit_freq_divider_1.dff_nclk_0.nCLK a_62654_21971# 0.31887f
C19 a_61394_23732# VDD 0.38531f
C20 charge_pump_0.vout VDD 0.06128f
C21 3bit_freq_divider_0.dff_nclk_0.nCLK a_54504_22015# 0.37259f
C22 a_53899_22244# VDD 0.26052f
C23 a_53022_43738# a_53058_43159# 0.24146f
C24 a_51693_23426# X1 0.01735f
C25 a_53065_23691# 3bit_freq_divider_0.dff_nclk_0.nCLK 0.29533f
C26 3bit_freq_divider_1.dff_nclk_0.nCLK 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.nQ 0.0874f
C27 3bit_freq_divider_0.EN a_59097_54704# 0.03561f
C28 a_57111_40283# VDD 1.36202f
C29 a_64383_23889# VDD 0.41974f
C30 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.Q a_54472_21129# 0.02559f
C31 a_61691_20534# a_62119_20605# 0.05314f
C32 a_51622_24863# 3bit_freq_divider_0.dff_nclk_0.nRST 0.10221f
C33 a_63463_23728# VDD 0.2349f
C34 a_51648_24041# a_51693_23075# 0.03957f
C35 a_62270_22299# VDD 0.26052f
C36 vco_wob_0.vctl a_53285_42591# 0.08086f
C37 a_53058_43159# a_53152_43159# 0.42803f
C38 a_53022_43738# a_54494_43159# 0.04f
C39 VDD CLK_OUT 0.38178f
C40 a_64384_21091# a_64714_21414# 0.014f
C41 m2_16847_2260# m3_16847_2260# 0.2063p
C42 a_53445_23726# VDD 0.31261f
C43 a_61887_20534# a_62900_20179# 0.04306f
C44 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.Q a_52886_21392# 0.12248f
C45 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.nQ a_53445_21970# 0.10118f
C46 a_53152_43159# a_54494_43159# 0.77984f
C47 a_58426_43159# a_57178_43159# 0.1057f
C48 vco_wob_0.vctl a_55770_40850# 0.05041f
C49 a_54504_23771# VDD 0.38531f
C50 a_53774_21934# 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.33731f
C51 3bit_freq_divider_0.freq_div_cell_0.Cin a_54472_22885# 0.01011f
C52 m5_17331_2744# m6_17427_2840# 84.0579f
C53 vco_wob_0.vctl a_57173_40413# 0.03129f
C54 a_51600_24907# a_51759_25014# 0.01952f
C55 m7_16847_2260# CLK_IN 1.44946f
C56 3bit_freq_divider_1.freq_div_cell_1.Cout a_61707_21488# 0.01154f
C57 a_51693_23426# a_51684_22284# 0.45825f
C58 a_51684_22692# X1 0.03873f
C59 a_63255_21488# Y2 0.39947f
C60 a_53968_20434# VDD 0.2982f
C61 a_53058_43159# VDD 1.37421f
C62 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.Q 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.D 0.22983f
C63 a_61887_20534# VDD 0.19386f
C64 a_51648_24041# a_51631_22774# 0.02302f
C65 a_61707_21488# a_61675_21130# 0.0104f
C66 3bit_freq_divider_0.freq_div_cell_0.Cout 3bit_freq_divider_0.freq_div_cell_1.Cout 0.09134f
C67 a_54494_43159# VDD 1.29885f
C68 VDD Y0 0.55412f
C69 3bit_freq_divider_0.dff_nclk_0.nCLK X2 0.64366f
C70 a_51759_25014# VDD 0.0834f
C71 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.D 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.40308f
C72 3bit_freq_divider_1.dff_nclk_0.nRST a_64419_23326# 0.16457f
C73 a_64383_23434# a_64419_23326# 0.66077f
C74 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.D a_61691_22290# 0.01446f
C75 a_51684_22692# a_51684_22284# 0.47248f
C76 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.Q a_63426_22886# 0.01011f
C77 m3_17285_2698# CLK_OUT 0.2919f
C78 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.Q Y2 0.15836f
C79 a_47777_29803# CLK_IN 0.17902f
C80 a_51631_22774# 3bit_freq_divider_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.33833f
C81 3bit_freq_divider_1.sg13g2_or3_1_0.C 3bit_freq_divider_1.dff_nclk_0.nCLK 0.13894f
C82 3bit_freq_divider_0.sg13g2_or3_1_0.B X2 0.33008f
C83 3bit_freq_divider_1.freq_div_cell_0.Cout a_61707_23244# 0.01154f
C84 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.sg13g2_dfrbp_1_0.CLK a_61394_23732# 0.08213f
C85 a_54434_24904# VDD 0.27564f
C86 vco_wob_0.vctl a_57178_43159# 0.026f
C87 charge_pump_0.bias_p a_58536_54976# 0.38944f
C88 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.Q Y1 0.18013f
C89 charge_pump_0.bias_n a_59097_54704# 0.01331f
C90 a_57112_40850# a_55831_40413# 0.23035f
C91 a_55862_56737# VDD 0.47223f
C92 a_61707_21488# 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.D 0.24715f
C93 a_56742_53480# a_56828_53480# 0.09853f
C94 a_54489_40413# a_53085_40283# 0.01232f
C95 a_53147_40413# a_54427_40283# 0.42019f
C96 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.Q a_52924_22885# 0.01011f
C97 a_53738_22270# a_54504_22015# 0.47248f
C98 a_53968_22190# a_53899_22244# 0.70262f
C99 a_63426_22886# VDD 0.20834f
C100 3bit_freq_divider_0.sg13g2_or3_1_0.A X2 0.2051f
C101 VDD X0 1.32697f
C102 3bit_freq_divider_0.dff_nclk_0.nCLK a_53065_21935# 0.31904f
C103 3bit_freq_divider_0.sg13g2_or3_1_0.C a_51648_21103# 0.25034f
C104 PFD_0.VCO_CLK a_46817_27899# 0.92547f
C105 a_48909_28913# a_47954_28913# 0.39061f
C106 a_61394_23732# a_62119_24117# 0.45825f
C107 a_58515_40413# a_58453_40283# 0.10827f
C108 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.Q a_52950_23913# 0.12519f
C109 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.D 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.40308f
C110 3bit_freq_divider_0.sg13g2_nand2_1_0.Y VDD 3.38843f
C111 m3_17285_2698# Y0 0.2919f
C112 a_61691_22290# a_62119_22361# 0.05314f
C113 a_56038_24617# VDD 0.0448f
C114 3bit_freq_divider_1.freq_div_cell_0.Cin 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.D 0.084f
C115 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.nQ a_53445_23726# 0.10118f
C116 a_53774_23690# a_53738_24026# 0.44698f
C117 a_61887_22290# a_62900_21935# 0.04306f
C118 3bit_freq_divider_0.dff_nclk_0.nCLK 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.D 0.21745f
C119 3bit_freq_divider_0.dff_nclk_0.nCLK a_52886_21392# 0.10313f
C120 3bit_freq_divider_1.dff_nclk_0.nCLK a_63426_21130# 0.03449f
C121 a_52950_22157# 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.nQ 0.21609f
C122 3bit_freq_divider_1.dff_nclk_0.nCLK 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.D 0.21745f
C123 a_53774_23690# 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.33731f
C124 a_53738_24026# a_53968_23946# 0.13068f
C125 a_64383_23628# VDD 0.62587f
C126 3bit_freq_divider_1.sg13g2_or3_1_0.C a_63426_24642# 0.10662f
C127 a_54494_43159# a_55969_42591# 0.03153f
C128 a_53022_43738# a_59800_40852# 0.01439f
C129 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.sg13g2_dfrbp_1_0.CLK VDD 0.27798f
C130 a_51622_24863# VDD 0.09559f
C131 a_64384_21091# VDD 0.34084f
C132 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.Q a_54472_24641# 0.02559f
C133 a_52944_43077# a_53147_40413# 0.40206f
C134 a_53022_43738# a_54427_40283# 0.18981f
C135 3bit_freq_divider_0.dff_nclk_0.nCLK X1 0.26228f
C136 a_53774_20178# VDD 0.67672f
C137 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.Q 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.D 0.22983f
C138 3bit_freq_divider_1.sg13g2_tiehi_1.L_HI a_60584_24580# 0.12404f
C139 3bit_freq_divider_0.dff_nclk_0.D a_51685_23725# 0.12409f
C140 3bit_freq_divider_0.dff_nclk_0.nCLK 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.D 0.21745f
C141 3bit_freq_divider_1.sg13g2_nand2_1_0.Y a_60967_23234# 0.08797f
C142 3bit_freq_divider_0.sg13g2_or3_1_0.C 3bit_freq_divider_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.28129f
C143 a_61707_23244# a_61878_22886# 0.36535f
C144 3bit_freq_divider_0.sg13g2_tiehi_1.L_HI VDD 0.77158f
C145 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.Q 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.nQ 0.02712f
C146 m3_17285_2698# X0 0.30224f
C147 a_61707_25000# VDD 0.27566f
C148 a_55941_24882# VDD 0.10494f
C149 a_63255_21488# a_63223_21130# 0.0104f
C150 3bit_freq_divider_1.sg13g2_or3_1_0.A a_64384_21091# 0.31317f
C151 3bit_freq_divider_0.sg13g2_or3_1_0.B X1 0.27832f
C152 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.Q 3bit_freq_divider_1.freq_div_cell_0.Cout 0.22232f
C153 a_64731_24890# 3bit_freq_divider_1.dff_nclk_0.nRST 0.01267f
C154 a_52886_21392# 3bit_freq_divider_0.sg13g2_or3_1_0.A 0.23182f
C155 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.Q a_63463_23728# 0.12519f
C156 3bit_freq_divider_0.dff_nclk_0.nRST a_51693_23075# 0.16442f
C157 3bit_freq_divider_1.dff_nclk_0.nCLK a_62900_23691# 0.24211f
C158 3bit_freq_divider_1.dff_nclk_0.nCLK a_62119_22361# 0.32758f
C159 a_63255_23244# Y2 0.01433f
C160 3bit_freq_divider_0.dff_nclk_0.nCLK a_53899_22244# 0.17328f
C161 a_64419_23326# a_64383_23300# 0.70262f
C162 charge_pump_0.vout a_56695_49467# 0.02916f
C163 a_54427_40283# VDD 1.36925f
C164 3bit_freq_divider_0.EN a_58734_56203# 0.07729f
C165 a_61691_20534# a_61887_20534# 0.45047f
C166 a_51648_24438# 3bit_freq_divider_0.dff_nclk_0.D 0.2233f
C167 a_64383_23889# 3bit_freq_divider_1.dff_nclk_0.D 0.09445f
C168 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.Q 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.D 0.22983f
C169 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.D a_53774_23690# 0.01446f
C170 m1_17285_2698# m2_17285_2698# 0.20496p
C171 a_53022_43738# a_52944_43077# 0.93638f
C172 3bit_freq_divider_0.dff_nclk_0.nCLK a_53445_23726# 0.24213f
C173 a_47777_29803# VDD 1.07957f
C174 3bit_freq_divider_1.dff_nclk_0.D CLK_OUT 0.01884f
C175 a_61887_20534# a_62654_20215# 0.40027f
C176 a_54434_24904# 3bit_freq_divider_0.freq_div_cell_0.Cin 0.01154f
C177 a_53065_21935# a_53738_22270# 0.40027f
C178 a_53774_21934# a_53445_21970# 0.04324f
C179 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.D a_61878_24642# 0.12185f
C180 a_62900_21935# VDD 0.30801f
C181 vco_wob_0.vctl a_53086_40850# 0.04284f
C182 a_52944_43077# a_53152_43159# 0.3548f
C183 a_57084_43159# a_55836_43159# 0.09926f
C184 3bit_freq_divider_0.dff_nclk_0.nCLK a_54504_23771# 0.37259f
C185 a_53899_24000# VDD 0.26493f
C186 3bit_freq_divider_1.freq_div_cell_0.Cout VDD 1.22849f
C187 3bit_freq_divider_1.sg13g2_or3_1_0.C a_64419_23326# 0.01089f
C188 vco_wob_0.vctl a_54489_40413# 0.04184f
C189 a_53065_20179# a_53774_20178# 0.02335f
C190 a_52950_20401# 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.nQ 0.21609f
C191 m5_16847_2260# m6_16847_2260# 0.13106p
C192 charge_pump_0.vout vco_wob_0.vctl 0.05724f
C193 m6_17427_2840# CLK_IN 1.23795f
C194 Y1 Y2 2.64011f
C195 3bit_freq_divider_1.dff_nclk_0.nCLK a_62270_20543# 0.17248f
C196 3bit_freq_divider_0.dff_nclk_0.nRST a_51631_22774# 0.3267f
C197 3bit_freq_divider_1.freq_div_cell_0.Cout 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.01369f
C198 3bit_freq_divider_0.dff_nclk_0.nCLK a_53968_20434# 0.32507f
C199 3bit_freq_divider_0.dff_nclk_0.D X1 0.11556f
C200 a_53738_20514# VDD 0.19386f
C201 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.Q Y0 0.20944f
C202 3bit_freq_divider_0.freq_div_cell_0.Cin 3bit_freq_divider_0.sg13g2_nand2_1_0.Y 0.25573f
C203 a_61394_20220# VDD 0.36995f
C204 PFD_0.DOWN a_54747_49259# 0.01456f
C205 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.D a_54504_22015# 0.3562f
C206 3bit_freq_divider_1.freq_div_cell_0.Cout a_60967_21478# 0.13034f
C207 a_52924_22885# VDD 0.20953f
C208 3bit_freq_divider_1.dff_nclk_0.nRST a_64384_24445# 0.04054f
C209 a_52944_43077# VDD 0.7984f
C210 3bit_freq_divider_0.EN 3bit_freq_divider_1.sg13g2_nand2_1_0.Y 0.12799f
C211 a_63463_20216# VDD 0.2331f
C212 a_52886_24904# VDD 0.28115f
C213 a_64398_24796# CLK_OUT 0.02652f
C214 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.Q a_61878_22886# 0.02559f
C215 3bit_freq_divider_0.EN X2 0.11756f
C216 3bit_freq_divider_0.dff_nclk_0.D a_51684_22284# 0.43097f
C217 3bit_freq_divider_0.sg13g2_nand2_1_0.Y 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.10521f
C218 a_45579_29803# CLK_IN 1.21724f
C219 3bit_freq_divider_1.sg13g2_or3_1_0.B VDD 0.10974f
C220 3bit_freq_divider_1.freq_div_cell_0.Cout a_61878_21130# 0.01011f
C221 vco_wob_0.vctl a_54494_43159# 0.0248f
C222 a_55770_40850# a_54489_40413# 0.23444f
C223 3bit_freq_divider_0.sg13g2_tiehi_1.L_HI 3bit_freq_divider_0.freq_div_cell_0.Cin 0.14552f
C224 a_63255_23244# Y1 0.39563f
C225 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.sg13g2_dfrbp_1_0.CLK a_61691_20534# 0.33731f
C226 a_53738_22270# a_53899_22244# 0.66077f
C227 a_54434_23148# 3bit_freq_divider_0.freq_div_cell_0.Cout 0.01154f
C228 3bit_freq_divider_1.dff_nclk_0.sg13g2_dfrbp_1_0.CLK VDD 0.28742f
C229 a_53065_20179# a_53738_20514# 0.40027f
C230 a_53774_20178# a_53445_20214# 0.04324f
C231 a_63255_25000# 3bit_freq_divider_1.sg13g2_or3_1_0.C 0.23357f
C232 3bit_freq_divider_1.sg13g2_or3_1_0.B 3bit_freq_divider_1.sg13g2_or3_1_0.A 0.72102f
C233 a_61878_22886# VDD 0.21321f
C234 a_52886_21392# X2 0.39847f
C235 a_57173_40413# a_57111_40283# 0.11922f
C236 a_61691_24046# a_62270_24055# 0.04304f
C237 a_61394_23732# a_61887_24046# 0.47248f
C238 a_53774_20178# 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.33731f
C239 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.Q 3bit_freq_divider_0.freq_div_cell_0.Cout 0.22232f
C240 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.nQ VDD 0.18275f
C241 3bit_freq_divider_0.dff_nclk_0.nCLK 3bit_freq_divider_0.sg13g2_nand2_1_0.Y 0.23907f
C242 a_62270_24055# a_62654_23727# 0.03957f
C243 a_52886_23148# a_53350_22885# 0.0104f
C244 a_61691_22290# a_61887_22290# 0.45047f
C245 3bit_freq_divider_0.sg13g2_or3_1_0.C 3bit_freq_divider_0.dff_nclk_0.nRST 0.57774f
C246 3bit_freq_divider_1.freq_div_cell_0.Cin a_61707_25000# 0.01154f
C247 a_53065_23691# a_53445_23726# 0.41048f
C248 3bit_freq_divider_1.freq_div_cell_1.Cout VDD 0.4595f
C249 a_61887_22290# a_62654_21971# 0.40027f
C250 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.D 3bit_freq_divider_1.sg13g2_nand2_1_0.Y 0.04726f
C251 a_46749_30782# a_47777_29803# 0.4544f
C252 a_45579_29803# a_45451_28860# 0.44406f
C253 X1 X2 0.01072f
C254 a_64459_24995# VDD 0.08543f
C255 a_51693_23075# VDD 0.2446f
C256 3bit_freq_divider_0.freq_div_cell_0.Cout a_54434_21392# 0.12082f
C257 3bit_freq_divider_1.dff_nclk_0.nRST VDD 0.60883f
C258 charge_pump_0.bias_p nEN 0.0229f
C259 a_64383_23434# VDD 0.19308f
C260 a_63255_25000# a_63426_24642# 0.36535f
C261 a_53152_43159# a_54627_42591# 0.03153f
C262 3bit_freq_divider_1.dff_nclk_0.D a_64383_23628# 0.03728f
C263 a_53738_24026# 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.01324f
C264 a_54434_23148# a_54898_22885# 0.0104f
C265 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.D a_54472_22885# 0.12185f
C266 3bit_freq_divider_0.CLK_IN a_58653_42591# 0.2448f
C267 a_53022_43738# a_58515_40413# 0.06975f
C268 3bit_freq_divider_0.dff_nclk_0.nCLK a_53774_20178# 0.35517f
C269 a_64383_23628# a_64424_22200# 0.17766f
C270 a_52950_20401# VDD 0.2331f
C271 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.Q a_61707_25000# 0.46099f
C272 a_60967_21478# 3bit_freq_divider_1.freq_div_cell_1.Cout 0.13166f
C273 a_60385_24717# a_60385_24947# 0.10864f
C274 a_54434_21392# 3bit_freq_divider_0.freq_div_cell_1.Cout 0.01154f
C275 a_52944_43077# a_53085_40283# 0.45412f
C276 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.Q a_52886_23148# 0.12248f
C277 3bit_freq_divider_0.EN X1 0.5347f
C278 3bit_freq_divider_1.freq_div_cell_0.Cin 3bit_freq_divider_1.freq_div_cell_0.Cout 0.10559f
C279 a_64459_24995# a_64362_24865# 0.10864f
C280 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.Q a_62654_21971# 0.01984f
C281 a_52924_24641# VDD 0.21522f
C282 a_51631_22774# VDD 0.62631f
C283 a_51693_23075# a_51693_23426# 0.70262f
C284 3bit_freq_divider_0.EN 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.D 0.02119f
C285 3bit_freq_divider_1.dff_nclk_0.nCLK a_61691_24046# 0.35198f
C286 a_54627_42591# VDD 0.01623f
C287 Y0 Y2 0.0326f
C288 a_64362_24865# 3bit_freq_divider_1.dff_nclk_0.nRST 0.03098f
C289 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.Q 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.nQ 0.02712f
C290 a_53445_20214# a_53738_20514# 0.04306f
C291 3bit_freq_divider_0.dff_nclk_0.D X0 0.1238f
C292 a_46817_27899# VDD 1.02029f
C293 3bit_freq_divider_1.dff_nclk_0.nCLK a_61887_22290# 0.18493f
C294 3bit_freq_divider_1.dff_nclk_0.nCLK a_62654_23727# 0.29516f
C295 a_56013_24979# a_56137_24678# 0.10864f
C296 a_58536_54976# VDD 0.98046f
C297 a_53738_20514# 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.01324f
C298 PFD_0.UP a_54357_49278# 0.30851f
C299 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.D VDD 0.9437f
C300 3bit_freq_divider_1.dff_nclk_0.nCLK 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.nQ 0.02503f
C301 a_54434_21392# a_54898_21129# 0.0104f
C302 a_58515_40413# VDD 1.36426f
C303 a_55948_56737# charge_pump_0.bias_p 0.02673f
C304 3bit_freq_divider_0.EN charge_pump_0.bias_n 0.02661f
C305 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.D a_54472_21129# 0.12185f
C306 a_61691_20534# a_61394_20220# 0.17766f
C307 a_51648_21103# a_51708_21413# 0.014f
C308 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK VDD 0.29872f
C309 a_61691_22290# VDD 0.68813f
C310 a_62270_24055# VDD 0.26494f
C311 a_53022_43738# a_57084_43159# 0.19696f
C312 m1_16847_2260# m2_16847_2260# 0.2063p
C313 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.Q VDD 1.68952f
C314 a_53774_23690# VDD 0.70098f
C315 a_45579_29803# VDD 0.45874f
C316 a_61887_20534# a_62119_20605# 0.13068f
C317 a_51684_22692# a_51693_23075# 0.66077f
C318 a_61707_25000# a_61878_24642# 0.36535f
C319 a_62654_21971# VDD 0.4336f
C320 a_64384_21091# a_64714_21300# 0.02055f
C321 a_55345_24897# VDD 0.45478f
C322 a_55742_43159# a_54494_43159# 0.10275f
C323 vco_wob_0.vctl a_57311_42591# 0.08436f
C324 a_53022_43738# 3bit_freq_divider_0.CLK_IN 0.16863f
C325 a_61707_23244# 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.D 0.24715f
C326 3bit_freq_divider_0.dff_nclk_0.nCLK a_53899_24000# 0.17312f
C327 a_53968_23946# VDD 0.32286f
C328 a_51631_22774# a_51693_23426# 0.05331f
C329 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK a_61691_22290# 0.33731f
C330 a_62654_20215# a_63463_20216# 0.09575f
C331 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.nQ VDD 0.18067f
C332 a_53065_21935# a_53899_22244# 0.03957f
C333 a_52950_20401# a_53065_20179# 0.09575f
C334 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.D 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.40308f
C335 vco_wob_0.vctl a_59800_40852# 0.05123f
C336 m4_17285_2698# m5_17331_2744# 0.1814p
C337 3bit_freq_divider_0.dff_nclk_0.nRST a_51648_24041# 0.30513f
C338 charge_pump_0.vout a_54357_49278# 0.01432f
C339 a_63463_20216# 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.nQ 0.21609f
C340 a_63463_23728# Y1 0.03561f
C341 m5_17331_2744# CLK_IN 0.42278f
C342 CLK_OUT Y1 0.01478f
C343 m6_16847_2260# m7_16847_2260# 39.787f
C344 3bit_freq_divider_1.dff_nclk_0.nCLK 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.Q 1.03922f
C345 3bit_freq_divider_0.dff_nclk_0.nCLK a_53738_20514# 0.18358f
C346 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.Q a_52950_20401# 0.12389f
C347 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.D a_54472_24641# 0.12185f
C348 a_54434_24904# a_54898_24641# 0.0104f
C349 3bit_freq_divider_1.dff_nclk_0.nCLK a_62900_20179# 0.2629f
C350 a_54504_20259# VDD 0.36995f
C351 3bit_freq_divider_0.dff_nclk_0.nCLK a_52924_22885# 0.03415f
C352 a_57084_43159# VDD 1.35049f
C353 a_51684_22692# a_51631_22774# 0.45006f
C354 3bit_freq_divider_0.dff_nclk_0.nRST 3bit_freq_divider_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.16209f
C355 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.D a_61878_21130# 0.12185f
C356 3bit_freq_divider_0.freq_div_cell_0.Cout VDD 1.22849f
C357 3bit_freq_divider_1.freq_div_cell_0.Cin a_61878_22886# 0.01011f
C358 3bit_freq_divider_0.CLK_IN VDD 1.60757f
C359 3bit_freq_divider_0.sg13g2_or3_1_0.C VDD 0.20391f
C360 a_51684_22284# X1 0.0269f
C361 3bit_freq_divider_0.sg13g2_or3_1_0.B a_52924_22885# 0.10697f
C362 a_60584_24580# VDD 0.10495f
C363 PFD_0.VCO_CLK 3bit_freq_divider_0.dff_nclk_0.nRST 0.06912f
C364 3bit_freq_divider_1.dff_nclk_0.nCLK VDD 2.89514f
C365 a_64383_23300# VDD 0.29403f
C366 Y0 Y1 1.97044f
C367 a_46817_27899# a_47954_28913# 0.22374f
C368 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.D a_61394_23732# 0.3562f
C369 3bit_freq_divider_1.freq_div_cell_0.Cout 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.Q 0.42266f
C370 3bit_freq_divider_0.sg13g2_nand2_1_0.Y a_55345_23141# 0.08797f
C371 3bit_freq_divider_1.dff_nclk_0.nCLK 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.60301f
C372 3bit_freq_divider_0.freq_div_cell_1.Cout VDD 0.4595f
C373 a_54428_40850# a_53147_40413# 0.23834f
C374 a_63255_23244# a_63426_22886# 0.36535f
C375 charge_pump_0.bias_n charge_pump_0.vout 0.23558f
C376 3bit_freq_divider_1.sg13g2_or3_1_0.C VDD 0.19202f
C377 a_58454_40850# a_58515_40413# 0.03243f
C378 3bit_freq_divider_1.sg13g2_nand2_1_0.Y 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.10521f
C379 3bit_freq_divider_1.dff_nclk_0.nCLK 3bit_freq_divider_1.sg13g2_or3_1_0.A 0.48568f
C380 a_51685_23725# X0 0.02143f
C381 3bit_freq_divider_1.dff_nclk_0.D 3bit_freq_divider_1.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.17618f
C382 a_52886_23148# VDD 0.25998f
C383 a_55831_40413# a_55769_40283# 0.12854f
C384 3bit_freq_divider_0.dff_nclk_0.nCLK 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.nQ 0.08742f
C385 a_64424_22200# 3bit_freq_divider_1.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.0838f
C386 a_53774_21934# VDD 0.69275f
C387 3bit_freq_divider_0.sg13g2_nand2_1_0.Y a_55345_21385# 0.08797f
C388 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.Q 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.D 0.22983f
C389 a_61691_22290# a_61394_21976# 0.17766f
C390 a_62270_24055# a_62119_24117# 0.70262f
C391 a_61691_24046# a_62900_23691# 0.04324f
C392 3bit_freq_divider_0.EN X0 0.11772f
C393 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.Q a_63463_20216# 0.12389f
C394 vco_wob_0.vctl a_60528_49446# 0.01545f
C395 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.Q 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.nQ 0.02712f
C396 3bit_freq_divider_1.sg13g2_tiehi_1.L_HI a_60967_24990# 0.21784f
C397 a_62654_23727# a_62900_23691# 0.41048f
C398 a_61887_22290# a_62119_22361# 0.13068f
C399 a_45579_29803# a_46749_30782# 0.25388f
C400 a_64383_23706# VDD 0.30655f
C401 3bit_freq_divider_0.EN 3bit_freq_divider_0.sg13g2_nand2_1_0.Y 0.12847f
C402 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.Q 3bit_freq_divider_0.freq_div_cell_0.Cin 0.22232f
C403 a_63426_22886# Y1 0.01971f
C404 3bit_freq_divider_0.CLK_IN m6_60810_42209# 0.11742f
C405 a_62900_23691# 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.nQ 0.10118f
C406 a_53065_23691# a_53899_24000# 0.03957f
C407 a_62900_21935# Y2 0.0145f
C408 a_45451_28860# PFD_0.VCO_CLK 0.12714f
C409 a_62654_21971# a_63463_21972# 0.09575f
C410 a_63426_24642# VDD 0.20944f
C411 a_51648_21103# VDD 0.34051f
C412 a_55345_24897# 3bit_freq_divider_0.freq_div_cell_0.Cin 0.13167f
C413 3bit_freq_divider_0.freq_div_cell_0.Cout 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.Q 0.42266f
C414 3bit_freq_divider_0.sg13g2_or3_1_0.C a_51684_22692# 0.03556f
C415 a_52944_43077# a_53285_42591# 0.03491f
C416 3bit_freq_divider_1.dff_nclk_0.nRST 3bit_freq_divider_1.dff_nclk_0.D 0.7629f
C417 3bit_freq_divider_0.CLK_IN 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.Q 0.02001f
C418 3bit_freq_divider_1.dff_nclk_0.D a_64383_23434# 0.0175f
C419 a_63463_21972# 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.nQ 0.21609f
C420 a_51648_24438# X0 0.01187f
C421 a_60967_23234# 3bit_freq_divider_1.freq_div_cell_0.Cout 0.13167f
C422 a_56828_53480# nEN 0.06208f
C423 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.D a_61691_20534# 0.01446f
C424 a_57178_43159# a_57311_42591# 0.22378f
C425 a_53022_43738# a_55831_40413# 0.04637f
C426 3bit_freq_divider_1.dff_nclk_0.nRST a_64424_22200# 0.34882f
C427 3bit_freq_divider_0.dff_nclk_0.nCLK a_52950_20401# 0.05883f
C428 a_64383_23434# a_64424_22200# 0.47248f
C429 a_63426_21130# VDD 0.20953f
C430 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.D VDD 0.97883f
C431 a_52924_21129# VDD 0.20953f
C432 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 3bit_freq_divider_1.dff_nclk_0.nCLK 0.60301f
C433 a_53022_43738# a_58453_40283# 0.19288f
C434 3bit_freq_divider_0.CLK_IN a_58454_40850# 0.02056f
C435 3bit_freq_divider_0.sg13g2_nand2_1_0.Y 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.D 0.05125f
C436 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.Q a_52950_22157# 0.12389f
C437 m1_17285_2698# X0 0.01061f
C438 a_51648_24041# VDD 0.41893f
C439 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.Q 3bit_freq_divider_0.freq_div_cell_1.Cout 0.2223f
C440 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.D 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.40308f
C441 3bit_freq_divider_1.sg13g2_nand2_1_0.Y 3bit_freq_divider_1.freq_div_cell_0.Cout 0.3426f
C442 X0 X1 0.55463f
C443 a_64459_24995# a_64398_24796# 0.0229f
C444 3bit_freq_divider_1.sg13g2_tiehi_1.L_HI VDD 0.7718f
C445 3bit_freq_divider_1.sg13g2_or3_1_0.A a_63426_21130# 0.10614f
C446 3bit_freq_divider_0.freq_div_cell_0.Cin 3bit_freq_divider_0.freq_div_cell_0.Cout 0.10559f
C447 m7_16847_2260# Y1 1.40976f
C448 3bit_freq_divider_1.dff_nclk_0.nCLK a_61394_21976# 0.37259f
C449 a_54428_40850# VDD 0.01457f
C450 3bit_freq_divider_1.dff_nclk_0.nCLK a_62119_24117# 0.32742f
C451 a_64398_24796# 3bit_freq_divider_1.dff_nclk_0.nRST 0.10221f
C452 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.Q a_54434_23148# 0.46099f
C453 charge_pump_0.bias_p VDD 2.67087f
C454 a_53445_21970# VDD 0.30838f
C455 3bit_freq_divider_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK VDD 0.28742f
C456 3bit_freq_divider_0.sg13g2_nand2_1_0.Y 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.D 0.05067f
C457 a_61707_21488# VDD 0.2676f
C458 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.Q 3bit_freq_divider_1.freq_div_cell_1.Cout 0.2223f
C459 a_55831_40413# VDD 1.08631f
C460 a_55862_56737# charge_pump_0.bias_n 0.34812f
C461 3bit_freq_divider_1.dff_nclk_0.nCLK a_63463_21972# 0.05956f
C462 a_54504_20259# 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.08213f
C463 3bit_freq_divider_1.sg13g2_or3_1_0.B Y2 0.1586f
C464 3bit_freq_divider_0.dff_nclk_0.nCLK 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.60301f
C465 a_53022_43738# a_54400_43159# 0.19723f
C466 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.Q 3bit_freq_divider_0.dff_nclk_0.nCLK 0.08441f
C467 a_53774_23690# 3bit_freq_divider_0.dff_nclk_0.nCLK 0.35198f
C468 a_52950_23913# VDD 0.24052f
C469 a_58453_40283# VDD 1.38336f
C470 a_61394_20220# a_62119_20605# 0.45825f
C471 3bit_freq_divider_0.dff_nclk_0.D a_51693_23075# 0.01591f
C472 a_62900_23691# VDD 0.31029f
C473 a_62119_22361# VDD 0.31854f
C474 a_56013_24979# VDD 0.11379f
C475 a_54400_43159# a_53152_43159# 0.09188f
C476 a_53022_43738# a_55836_43159# 0.04103f
C477 vco_wob_0.vctl a_54627_42591# 0.07714f
C478 3bit_freq_divider_0.dff_nclk_0.nCLK a_53968_23946# 0.32517f
C479 PFD_0.VCO_CLK VDD 1.82327f
C480 a_53738_24026# VDD 0.22151f
C481 a_64419_23326# VDD 0.2446f
C482 PFD_0.DOWN PFD_0.VCO_CLK 0.20401f
C483 a_53774_21934# a_53968_22190# 0.05314f
C484 a_58426_43159# 3bit_freq_divider_0.CLK_IN 0.4131f
C485 vco_wob_0.vctl a_57112_40850# 0.05026f
C486 m4_16847_2260# m5_16847_2260# 0.2063p
C487 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.sg13g2_dfrbp_1_0.CLK VDD 0.30706f
C488 3bit_freq_divider_1.freq_div_cell_0.Cin 3bit_freq_divider_1.dff_nclk_0.nCLK 0.32366f
C489 m4_17285_2698# CLK_IN 0.39515f
C490 3bit_freq_divider_1.dff_nclk_0.nCLK a_61691_20534# 0.35517f
C491 vco_wob_0.vctl a_58515_40413# 0.02267f
C492 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.D a_53774_20178# 0.01446f
C493 3bit_freq_divider_1.dff_nclk_0.nCLK a_62654_20215# 0.31114f
C494 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.Q a_52924_21129# 0.01011f
C495 a_54472_24641# VDD 0.214f
C496 a_53899_20488# VDD 0.24492f
C497 VDD nEN 3.87548f
C498 3bit_freq_divider_0.dff_nclk_0.nCLK a_54504_20259# 0.37259f
C499 a_51648_24041# a_51684_22692# 0.40027f
C500 3bit_freq_divider_1.dff_nclk_0.nCLK 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.nQ 0.08552f
C501 a_54400_43159# VDD 1.37065f
C502 a_62270_20543# VDD 0.24492f
C503 3bit_freq_divider_0.dff_nclk_0.D a_51631_22774# 0.03728f
C504 a_61707_21488# a_61878_21130# 0.36535f
C505 3bit_freq_divider_0.dff_nclk_0.nCLK 3bit_freq_divider_0.freq_div_cell_0.Cout 0.32366f
C506 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.Q 3bit_freq_divider_1.dff_nclk_0.nCLK 0.0844f
C507 a_55836_43159# VDD 1.00781f
C508 a_64383_23889# a_64383_23628# 0.02302f
C509 a_61707_25000# 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.D 0.24715f
C510 3bit_freq_divider_0.sg13g2_or3_1_0.C 3bit_freq_divider_0.dff_nclk_0.nCLK 0.13894f
C511 a_63255_23244# 3bit_freq_divider_1.sg13g2_or3_1_0.B 0.23215f
C512 a_51721_24988# VDD 0.08543f
C513 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.Q 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.D 0.22983f
C514 a_56137_24678# VDD 0.11858f
C515 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.D a_61394_21976# 0.3562f
C516 a_51684_22692# 3bit_freq_divider_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.01473f
C517 3bit_freq_divider_1.dff_nclk_0.nCLK 3bit_freq_divider_1.dff_nclk_0.D 0.04354f
C518 3bit_freq_divider_1.dff_nclk_0.D a_64383_23300# 0.04146f
C519 a_62654_21971# 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.Q 0.0119f
C520 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.Q 3bit_freq_divider_1.sg13g2_or3_1_0.C 0.05745f
C521 a_45451_28860# CLK_IN 0.13923f
C522 3bit_freq_divider_1.sg13g2_nand2_1_0.Y 3bit_freq_divider_1.freq_div_cell_1.Cout 0.07626f
C523 a_45658_27900# a_46817_27899# 0.43194f
C524 m7_16847_2260# CLK_OUT 1.40976f
C525 3bit_freq_divider_0.sg13g2_or3_1_0.C 3bit_freq_divider_0.sg13g2_or3_1_0.B 1.00414f
C526 a_64383_23300# a_64424_22200# 0.45825f
C527 PFD_0.UP a_47777_29803# 0.62819f
C528 vco_wob_0.vctl 3bit_freq_divider_0.CLK_IN 0.50349f
C529 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.D VDD 0.97078f
C530 charge_pump_0.bias_n a_56742_53480# 0.05592f
C531 charge_pump_0.bias_p a_59097_54704# 0.04726f
C532 a_58734_56203# a_58536_54976# 0.19076f
C533 a_63255_25000# VDD 0.26507f
C534 a_57112_40850# a_57173_40413# 0.03159f
C535 3bit_freq_divider_1.sg13g2_or3_1_0.B Y1 0.13266f
C536 a_55948_56737# VDD 0.31573f
C537 3bit_freq_divider_1.dff_nclk_0.nCLK a_63255_21488# 0.10313f
C538 a_54489_40413# a_54427_40283# 0.12991f
C539 3bit_freq_divider_0.dff_nclk_0.nCLK a_52886_23148# 0.10223f
C540 a_57173_40413# a_58515_40413# 0.58365f
C541 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.sg13g2_dfrbp_1_0.CLK a_61887_20534# 0.01324f
C542 a_53738_22270# 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.01324f
C543 a_53774_20178# a_53968_20434# 0.05314f
C544 a_53065_20179# a_53899_20488# 0.03957f
C545 3bit_freq_divider_0.dff_nclk_0.nCLK a_53774_21934# 0.35569f
C546 a_52950_22157# VDD 0.2364f
C547 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.Q a_61707_23244# 0.46099f
C548 PFD_0.VCO_CLK a_47954_28913# 1.24436f
C549 a_61887_24046# a_62270_24055# 0.66077f
C550 a_61691_24046# a_62654_23727# 0.02302f
C551 a_58515_40413# a_59799_40285# 0.46077f
C552 a_51759_25014# a_51622_24863# 0.14868f
C553 a_51600_24907# 3bit_freq_divider_0.dff_nclk_0.nRST 0.01267f
C554 a_54504_22015# 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.08213f
C555 a_54842_49733# VDD 0.03367f
C556 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.Q a_63426_24642# 0.02246f
C557 a_52924_22885# X1 0.02265f
C558 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.Q a_53065_23691# 0.02071f
C559 a_56887_49467# a_56695_49467# 0.01287f
C560 a_61394_21976# a_62119_22361# 0.45825f
C561 a_53065_23691# a_53774_23690# 0.02335f
C562 a_52950_23913# 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.nQ 0.21609f
C563 a_60385_24558# VDD 0.04481f
C564 3bit_freq_divider_0.CLK_IN 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.Q 0.02001f
C565 a_52886_23148# 3bit_freq_divider_0.sg13g2_or3_1_0.B 0.23215f
C566 3bit_freq_divider_1.dff_nclk_0.D a_64383_23706# 0.12409f
C567 3bit_freq_divider_1.sg13g2_tiehi_1.L_HI 3bit_freq_divider_1.freq_div_cell_0.Cin 0.14552f
C568 m7_16847_2260# Y0 1.40976f
C569 a_62654_23727# 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.nQ 0.05822f
C570 a_54434_23148# VDD 0.2676f
C571 a_64731_24890# VDD 0.04155f
C572 3bit_freq_divider_0.dff_nclk_0.nCLK a_51648_21103# 0.33244f
C573 a_62654_21971# Y2 0.02368f
C574 3bit_freq_divider_0.EN 3bit_freq_divider_1.freq_div_cell_1.Cout 0.01552f
C575 a_53065_21935# 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.nQ 0.0571f
C576 3bit_freq_divider_1.dff_nclk_0.nCLK 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.Q 1.04018f
C577 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.nQ Y2 0.04365f
C578 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.Q VDD 1.42273f
C579 a_53022_43738# a_53147_40413# 0.08011f
C580 3bit_freq_divider_0.dff_nclk_0.nRST VDD 0.60215f
C581 3bit_freq_divider_0.freq_div_cell_0.Cin 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.01369f
C582 a_55836_43159# a_55969_42591# 0.22378f
C583 a_52944_43077# a_53086_40850# 0.23665f
C584 3bit_freq_divider_1.sg13g2_nand2_1_0.Y 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.D 0.05067f
C585 a_61707_23244# VDD 0.2676f
C586 charge_pump_0.vout a_54747_49259# 0.13589f
C587 3bit_freq_divider_0.dff_nclk_0.nCLK a_52924_21129# 0.03449f
C588 a_53022_43738# a_55769_40283# 0.19098f
C589 3bit_freq_divider_0.sg13g2_or3_1_0.B a_51648_21103# 0.26158f
C590 VDD CLK_IN 2.49441f
C591 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.nQ VDD 0.18065f
C592 3bit_freq_divider_1.sg13g2_tiehi_1.L_HI 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.Q 0.42892f
C593 a_54434_21392# VDD 0.2676f
C594 PFD_0.DOWN CLK_IN 0.06328f
C595 3bit_freq_divider_0.sg13g2_tiehi_1.L_HI a_54434_24904# 0.12082f
C596 a_51685_23725# a_51631_22774# 0.04324f
C597 a_62654_23727# 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.Q 0.0119f
C598 a_64362_24865# a_64731_24890# 0.01952f
C599 3bit_freq_divider_0.CLK_IN a_59799_40285# 0.11621f
C600 a_60479_25023# VDD 0.01215f
C601 a_63255_21488# a_63426_21130# 0.36535f
C602 m7_16847_2260# X0 1.44946f
C603 m6_17427_2840# Y1 1.19758f
C604 3bit_freq_divider_1.dff_nclk_0.nCLK a_61887_24046# 0.18489f
C605 a_51648_21103# 3bit_freq_divider_0.sg13g2_or3_1_0.A 0.31317f
C606 a_53738_20514# a_53968_20434# 0.13068f
C607 3bit_freq_divider_0.dff_nclk_0.nCLK a_53445_21970# 0.27428f
C608 3bit_freq_divider_0.dff_nclk_0.nRST a_51693_23426# 0.3148f
C609 3bit_freq_divider_0.dff_nclk_0.nCLK 3bit_freq_divider_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.10701f
C610 a_53147_40413# VDD 0.81739f
C611 3bit_freq_divider_1.dff_nclk_0.nCLK Y2 0.86741f
C612 a_61691_24046# VDD 0.69635f
C613 charge_pump_0.vout a_60528_49446# 0.01545f
C614 a_55769_40283# VDD 1.37334f
C615 3bit_freq_divider_0.EN a_58536_54976# 0.21462f
C616 a_64384_24445# VDD 0.24105f
C617 a_51693_23075# X1 0.01284f
C618 a_61691_20534# a_62270_20543# 0.04304f
C619 a_61394_20220# a_61887_20534# 0.47248f
C620 a_52886_24904# a_53350_24641# 0.0104f
C621 3bit_freq_divider_0.sg13g2_or3_1_0.A a_52924_21129# 0.10614f
C622 a_61887_22290# VDD 0.21577f
C623 a_62654_23727# VDD 0.43765f
C624 3bit_freq_divider_0.EN 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.D 0.02092f
C625 a_53058_43159# a_52944_43077# 0.08875f
C626 a_53022_43738# a_53152_43159# 0.08218f
C627 3bit_freq_divider_0.dff_nclk_0.nCLK a_53738_24026# 0.18638f
C628 a_45451_28860# VDD 0.05543f
C629 3bit_freq_divider_0.CLK_IN 3bit_freq_divider_1.sg13g2_nand2_1_0.Y 0.2618f
C630 a_62270_20543# a_62654_20215# 0.03957f
C631 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.D 3bit_freq_divider_0.freq_div_cell_0.Cin 0.084f
C632 3bit_freq_divider_1.dff_nclk_0.D a_64419_23326# 0.01591f
C633 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.nQ VDD 0.18204f
C634 a_53774_21934# a_53738_22270# 0.44698f
C635 a_57084_43159# a_57178_43159# 0.42665f
C636 vco_wob_0.vctl a_54428_40850# 0.04894f
C637 m3_17285_2698# m4_17285_2698# 0.20496p
C638 3bit_freq_divider_1.sg13g2_tiehi_1.L_HI a_61878_24642# 0.01011f
C639 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.Q a_63426_21130# 0.01011f
C640 3bit_freq_divider_0.dff_nclk_0.nCLK 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.60301f
C641 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK a_61887_22290# 0.01324f
C642 m3_17285_2698# CLK_IN 0.30224f
C643 3bit_freq_divider_0.dff_nclk_0.nRST a_51684_22692# 0.126f
C644 a_55345_23141# 3bit_freq_divider_0.freq_div_cell_0.Cout 0.13167f
C645 3bit_freq_divider_1.sg13g2_nand2_1_0.Y 3bit_freq_divider_1.dff_nclk_0.nCLK 0.23907f
C646 a_53774_21934# a_54504_22015# 0.17766f
C647 a_53065_20179# 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.nQ 0.0571f
C648 a_57178_43159# 3bit_freq_divider_0.CLK_IN 0.20831f
C649 vco_wob_0.vctl a_55831_40413# 0.04109f
C650 3bit_freq_divider_1.dff_nclk_0.nCLK a_62119_20605# 0.32732f
C651 3bit_freq_divider_0.sg13g2_or3_1_0.C X2 0.04643f
C652 a_60967_24990# VDD 0.4548f
C653 3bit_freq_divider_0.dff_nclk_0.nCLK a_53899_20488# 0.17248f
C654 a_51648_24041# 3bit_freq_divider_0.dff_nclk_0.D 0.09445f
C655 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.Q 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.nQ 0.02712f
C656 a_53022_43738# VDD 13.1862f
C657 a_51631_22774# X1 0.02271f
C658 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.Q a_54434_21392# 0.46099f
C659 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.D 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.40308f
C660 a_60385_24947# a_60584_24580# 0.0229f
C661 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.Q VDD 1.41895f
C662 3bit_freq_divider_1.dff_nclk_0.nRST a_64383_23889# 0.30513f
C663 3bit_freq_divider_0.freq_div_cell_0.Cout a_55345_21385# 0.13034f
C664 a_53152_43159# VDD 1.05457f
C665 3bit_freq_divider_0.sg13g2_tiehi_1.L_HI a_55941_24882# 0.12404f
C666 a_64383_23889# a_64383_23434# 0.40027f
C667 a_62900_20179# VDD 0.30479f
C668 3bit_freq_divider_1.dff_nclk_0.nCLK a_63255_23244# 0.10223f
C669 a_51600_24907# VDD 0.04155f
C670 3bit_freq_divider_0.freq_div_cell_0.Cin a_54434_23148# 0.12082f
C671 3bit_freq_divider_1.dff_nclk_0.nRST CLK_OUT 0.07748f
C672 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.Q a_61707_21488# 0.46099f
C673 3bit_freq_divider_0.freq_div_cell_0.Cin 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.Q 0.42266f
C674 3bit_freq_divider_0.EN 3bit_freq_divider_0.CLK_IN 0.41907f
C675 3bit_freq_divider_0.dff_nclk_0.D 3bit_freq_divider_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.17618f
C676 a_63426_21130# Y2 0.02209f
C677 a_52886_24904# X0 0.40762f
C678 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.Q X1 0.01869f
C679 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.Q a_63255_25000# 0.14987f
C680 a_51631_22774# a_51684_22284# 0.17766f
C681 a_46749_30782# CLK_IN 0.97391f
C682 m6_17427_2840# CLK_OUT 1.19758f
C683 a_55345_21385# 3bit_freq_divider_0.freq_div_cell_1.Cout 0.13166f
C684 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.sg13g2_dfrbp_1_0.CLK a_61691_24046# 0.33731f
C685 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.D 3bit_freq_divider_0.dff_nclk_0.nCLK 0.21603f
C686 vco_wob_0.vctl a_55836_43159# 0.02497f
C687 charge_pump_0.bias_n a_58536_54976# 0.02549f
C688 charge_pump_0.bias_p a_58734_56203# 0.03822f
C689 PFD_0.VCO_CLK 3bit_freq_divider_0.dff_nclk_0.D 0.01884f
C690 3bit_freq_divider_0.freq_div_cell_0.Cout a_54472_21129# 0.01011f
C691 3bit_freq_divider_1.dff_nclk_0.nCLK Y1 0.23798f
C692 PFD_0.DOWN VDD 1.56226f
C693 a_55770_40850# a_55831_40413# 0.03778f
C694 a_53445_21970# a_53738_22270# 0.04306f
C695 3bit_freq_divider_0.EN 3bit_freq_divider_0.freq_div_cell_1.Cout 0.01552f
C696 3bit_freq_divider_1.sg13g2_or3_1_0.B a_63426_22886# 0.10697f
C697 a_55831_40413# a_57173_40413# 0.7336f
C698 a_53147_40413# a_53085_40283# 0.10818f
C699 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.sg13g2_dfrbp_1_0.CLK a_61394_20220# 0.08213f
C700 3bit_freq_divider_1.freq_div_cell_0.Cin a_61707_23244# 0.12082f
C701 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.D 3bit_freq_divider_0.freq_div_cell_0.Cout 0.084f
C702 a_53774_20178# a_53738_20514# 0.44698f
C703 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.nQ a_53445_20214# 0.10118f
C704 3bit_freq_divider_1.sg13g2_nand2_1_0.Y 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.D 0.05125f
C705 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK VDD 0.29872f
C706 3bit_freq_divider_0.dff_nclk_0.nCLK a_52950_22157# 0.05957f
C707 a_61691_24046# a_62119_24117# 0.05314f
C708 PFD_0.VCO_CLK a_45658_27900# 0.17296f
C709 a_57173_40413# a_58453_40283# 0.46167f
C710 3bit_freq_divider_1.sg13g2_or3_1_0.C Y1 0.16352f
C711 3bit_freq_divider_1.sg13g2_or3_1_0.A VDD 0.12797f
C712 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.D a_54504_20259# 0.3562f
C713 a_52950_23913# a_53065_23691# 0.09575f
C714 a_60967_21478# VDD 0.45855f
C715 a_61887_24046# a_62900_23691# 0.04306f
C716 a_61691_22290# a_62270_22299# 0.04304f
C717 a_61394_21976# a_61887_22290# 0.47248f
C718 a_52924_21129# X2 0.02265f
C719 a_62270_22299# a_62654_21971# 0.03957f
C720 m6_17427_2840# Y0 1.19758f
C721 a_53774_23690# a_53445_23726# 0.04324f
C722 a_53065_23691# a_53738_24026# 0.40027f
C723 a_64362_24865# VDD 0.08341f
C724 a_62900_23691# Y2 0.01917f
C725 3bit_freq_divider_0.sg13g2_or3_1_0.C X1 0.20623f
C726 a_51693_23426# VDD 0.29403f
C727 a_53065_21935# a_53774_21934# 0.02335f
C728 3bit_freq_divider_1.sg13g2_or3_1_0.B a_64384_21091# 0.26158f
C729 a_53774_23690# a_54504_23771# 0.17766f
C730 3bit_freq_divider_0.dff_nclk_0.nCLK 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.Q 1.03924f
C731 a_54494_43159# a_54627_42591# 0.22378f
C732 a_53968_23946# a_54504_23771# 0.45825f
C733 a_61878_21130# VDD 0.21321f
C734 a_53022_43738# a_53085_40283# 0.23019f
C735 a_64383_23628# 3bit_freq_divider_1.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.33833f
C736 a_53065_20179# VDD 0.42601f
C737 a_63426_24642# Y1 0.01474f
C738 3bit_freq_divider_0.dff_nclk_0.nCLK 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.nQ 0.08555f
C739 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.D a_53774_21934# 0.01446f
C740 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.D 3bit_freq_divider_1.dff_nclk_0.nCLK 0.21603f
C741 a_51648_24041# a_51685_23725# 0.41048f
C742 a_60385_24717# a_60584_24580# 0.14868f
C743 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.D 3bit_freq_divider_0.freq_div_cell_1.Cout 0.04623f
C744 m6_60810_42209# VDD 0.03757f
C745 a_51684_22692# VDD 0.19308f
C746 a_61707_23244# a_61675_22886# 0.0104f
C747 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.Q VDD 1.42261f
C748 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.Q a_63463_21972# 0.12389f
C749 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.sg13g2_dfrbp_1_0.CLK VDD 0.3071f
C750 a_52886_23148# X1 0.39847f
C751 m5_17331_2744# Y1 0.40842f
C752 m6_17427_2840# X0 1.23795f
C753 3bit_freq_divider_1.dff_nclk_0.nCLK a_61394_23732# 0.37259f
C754 a_55969_42591# VDD 0.0108f
C755 a_60967_24990# 3bit_freq_divider_1.freq_div_cell_0.Cin 0.13167f
C756 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.Q a_62654_23727# 0.02071f
C757 a_47954_28913# VDD 0.45155f
C758 a_52924_24641# X0 0.02265f
C759 3bit_freq_divider_1.dff_nclk_0.nCLK a_62270_22299# 0.17328f
C760 3bit_freq_divider_1.dff_nclk_0.nRST a_64383_23628# 0.3268f
C761 a_53968_20434# a_54504_20259# 0.45825f
C762 a_53968_22190# VDD 0.31854f
C763 a_64383_23434# a_64383_23628# 0.44985f
C764 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.Q 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.nQ 0.02712f
C765 a_53085_40283# VDD 1.35573f
C766 3bit_freq_divider_0.EN charge_pump_0.bias_p 0.33628f
C767 a_52886_21392# a_52924_21129# 0.36535f
C768 a_51648_24438# a_51648_24041# 0.09575f
C769 a_51648_21103# a_51708_21299# 0.02055f
C770 3bit_freq_divider_1.freq_div_cell_0.Cin 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.Q 0.42266f
C771 a_62119_24117# VDD 0.32287f
C772 a_64384_24445# 3bit_freq_divider_1.dff_nclk_0.D 0.2233f
C773 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.Q a_54434_24904# 0.46099f
C774 a_61394_21976# VDD 0.38024f
C775 a_53022_43738# a_58426_43159# 0.10045f
C776 a_46749_30782# VDD 1.12191f
C777 a_51684_22692# a_51693_23426# 0.13068f
C778 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.nQ VDD 0.18755f
C779 a_62270_20543# a_62119_20605# 0.70262f
C780 a_61691_20534# a_62900_20179# 0.04324f
C781 a_53065_21935# a_53445_21970# 0.41048f
C782 a_63463_21972# VDD 0.2345f
C783 3bit_freq_divider_0.freq_div_cell_0.Cin VDD 1.21627f
C784 a_55742_43159# a_55836_43159# 0.42148f
C785 m3_16847_2260# m4_16847_2260# 0.2063p
C786 vco_wob_0.vctl a_58653_42591# 0.08336f
C787 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.Q a_60967_24990# 0.30546f
C788 a_63255_25000# Y2 0.02709f
C789 charge_pump_0.bias_p a_54357_49278# 0.01013f
C790 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK a_61394_21976# 0.08213f
C791 a_62654_20215# a_62900_20179# 0.41048f
C792 a_53774_21934# a_53899_22244# 0.04304f
C793 a_55836_43159# a_57178_43159# 0.91818f
C794 vco_wob_0.vctl a_53147_40413# 0.04038f
C795 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.Q X0 0.24362f
C796 3bit_freq_divider_0.dff_nclk_0.nRST 3bit_freq_divider_0.dff_nclk_0.D 0.76289f
C797 a_62900_20179# 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.nQ 0.10118f
C798 charge_pump_0.vout a_56887_49467# 0.63953f
C799 3bit_freq_divider_1.dff_nclk_0.nCLK a_61887_20534# 0.18209f
C800 3bit_freq_divider_0.sg13g2_nand2_1_0.Y 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.11142f
C801 m6_17427_2840# m7_16847_2260# 25.5177f
C802 a_53445_20214# VDD 0.30479f
C803 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.Q a_53065_20179# 0.01984f
C804 3bit_freq_divider_1.freq_div_cell_0.Cin VDD 1.21632f
C805 a_64383_23889# a_64383_23706# 0.41048f
C806 a_61691_20534# VDD 0.67211f
C807 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.sg13g2_dfrbp_1_0.CLK VDD 0.27798f
C808 PFD_0.VCO_CLK a_51648_24438# 0.11636f
C809 a_58426_43159# VDD 1.36969f
C810 3bit_freq_divider_0.EN nEN 0.24728f
C811 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.D 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.40308f
C812 a_62654_20215# VDD 0.42601f
C813 3bit_freq_divider_1.freq_div_cell_0.Cout 3bit_freq_divider_1.freq_div_cell_1.Cout 0.09134f
C814 a_53065_23691# 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.Q 0.0119f
C815 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.nQ VDD 0.18065f
C816 3bit_freq_divider_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK X1 0.02018f
C817 a_60385_24717# 3bit_freq_divider_1.sg13g2_tiehi_1.L_HI 0.02161f
C818 3bit_freq_divider_1.sg13g2_or3_1_0.C Y0 0.12518f
C819 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.Q VDD 1.66358f
C820 vco_wob_0.vctl a_53022_43738# 0.09057f
C821 m5_17331_2744# CLK_OUT 0.40842f
C822 3bit_freq_divider_0.sg13g2_or3_1_0.C X0 0.41386f
C823 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.Q 3bit_freq_divider_0.sg13g2_tiehi_1.L_HI 0.42892f
C824 vco_wob_0.vctl a_53152_43159# 0.02282f
C825 3bit_freq_divider_0.dff_nclk_0.nCLK VDD 2.90191f
C826 3bit_freq_divider_0.sg13g2_nand2_1_0.Y 3bit_freq_divider_0.freq_div_cell_0.Cout 0.3426f
C827 3bit_freq_divider_0.CLK_IN 3bit_freq_divider_0.sg13g2_nand2_1_0.Y 0.2618f
C828 charge_pump_0.bias_n charge_pump_0.bias_p 1.09436f
C829 a_54428_40850# a_54489_40413# 0.03943f
C830 3bit_freq_divider_1.dff_nclk_0.nCLK a_63426_22886# 0.03415f
C831 3bit_freq_divider_1.dff_nclk_0.D VDD 0.84615f
C832 3bit_freq_divider_0.sg13g2_tiehi_1.L_HI a_55345_24897# 0.21784f
C833 charge_pump_0.bias_p charge_pump_0.vout 0.02402f
C834 a_51684_22284# 3bit_freq_divider_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.0838f
C835 a_59800_40852# a_58515_40413# 0.21632f
C836 a_54489_40413# a_55831_40413# 0.72984f
C837 a_64424_22200# VDD 0.36995f
C838 a_53065_20179# a_53445_20214# 0.41048f
C839 a_63426_24642# Y0 0.01851f
C840 a_55948_56737# 3bit_freq_divider_0.EN 0.0294f
C841 a_61691_24046# a_61887_24046# 0.45047f
C842 3bit_freq_divider_0.sg13g2_or3_1_0.B VDD 0.11082f
C843 a_55831_40413# a_57111_40283# 0.45955f
C844 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.Q a_55345_23141# 0.30546f
C845 a_53774_20178# a_54504_20259# 0.17766f
C846 a_63255_25000# Y1 0.01849f
C847 3bit_freq_divider_0.sg13g2_nand2_1_0.Y 3bit_freq_divider_0.freq_div_cell_1.Cout 0.07626f
C848 a_63255_21488# VDD 0.26051f
C849 a_61887_24046# a_62654_23727# 0.40027f
C850 vco_wob_0.vctl VDD 0.2823f
C851 m5_17331_2744# Y0 0.40842f
C852 3bit_freq_divider_1.freq_div_cell_0.Cin 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.01369f
C853 a_64383_23889# a_64419_23326# 0.03957f
C854 a_62270_22299# a_62119_22361# 0.70262f
C855 a_61691_22290# a_62900_21935# 0.04324f
C856 a_62654_23727# Y2 0.02178f
C857 a_61878_24642# VDD 0.21401f
C858 a_64383_23628# a_64383_23300# 0.05314f
C859 3bit_freq_divider_1.dff_nclk_0.nCLK 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.60301f
C860 a_52950_22157# a_53065_21935# 0.09575f
C861 3bit_freq_divider_1.dff_nclk_0.nCLK a_64384_21091# 0.33258f
C862 a_53022_43738# a_53285_42591# 0.02036f
C863 a_53445_23726# a_53738_24026# 0.04306f
C864 a_53774_23690# a_53899_24000# 0.04304f
C865 a_48909_28913# PFD_0.VCO_CLK 0.1514f
C866 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.nQ Y2 0.04535f
C867 a_62654_21971# a_62900_21935# 0.41048f
C868 3bit_freq_divider_0.sg13g2_or3_1_0.A VDD 0.12791f
C869 a_64398_24796# VDD 0.09559f
C870 charge_pump_0.bias_n nEN 0.06869f
C871 a_52886_24904# a_52924_24641# 0.36535f
C872 a_63255_25000# a_63223_24642# 0.0104f
C873 3bit_freq_divider_0.dff_nclk_0.nRST a_51685_23725# 0.25925f
C874 a_53152_43159# a_53285_42591# 0.22378f
C875 a_53738_24026# a_54504_23771# 0.47248f
C876 a_53968_23946# a_53899_24000# 0.70262f
C877 a_62900_21935# 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.nQ 0.10118f
C878 a_63255_21488# 3bit_freq_divider_1.sg13g2_or3_1_0.A 0.23182f
C879 a_54434_23148# a_54472_22885# 0.36535f
C880 a_53022_43738# a_57173_40413# 0.04406f
C881 a_57178_43159# a_58653_42591# 0.03205f
C882 3bit_freq_divider_1.dff_nclk_0.nRST 3bit_freq_divider_1.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.16234f
C883 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.D a_61394_20220# 0.3562f
C884 3bit_freq_divider_0.dff_nclk_0.nCLK a_53065_20179# 0.31132f
C885 a_64383_23434# 3bit_freq_divider_1.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.01473f
C886 a_54504_23771# 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.08213f
C887 a_64714_21300# VDD 0.01263f
C888 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.Q VDD 1.4225f
C889 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.Q a_54472_22885# 0.02559f
C890 3bit_freq_divider_1.sg13g2_or3_1_0.C a_64384_21091# 0.25034f
C891 3bit_freq_divider_0.CLK_IN a_59800_40852# 0.13041f
C892 a_53022_43738# a_59799_40285# 0.19389f
C893 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.Q a_53065_21935# 0.01984f
C894 3bit_freq_divider_0.dff_nclk_0.D VDD 0.84532f
C895 3bit_freq_divider_0.dff_nclk_0.nCLK 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.Q 1.0402f
C896 a_52886_21392# a_53350_21129# 0.0104f
C897 3bit_freq_divider_0.EN CLK_IN 0.09396f
C898 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.Q a_52886_24904# 0.14987f
C899 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.Q Y2 0.20327f
C900 m4_17285_2698# Y1 0.3817f
C901 m5_17331_2744# X0 0.42278f
C902 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.Q a_60967_23234# 0.30546f
C903 a_54434_23148# 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.D 0.24715f
C904 a_64362_24865# a_64398_24796# 0.14868f
C905 a_64383_23706# a_64383_23628# 0.04324f
C906 3bit_freq_divider_0.dff_nclk_0.nRST a_51648_24438# 0.04054f
C907 a_51648_24041# X0 0.0271f
C908 a_45658_27900# VDD 1.00659f
C909 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.Q a_60967_21478# 0.30546f
C910 a_55770_40850# VDD 0.01475f
C911 PFD_0.DOWN a_45658_27900# 0.61911f
C912 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.Q 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.D 0.22983f
C913 3bit_freq_divider_1.dff_nclk_0.nRST a_64383_23434# 0.126f
C914 a_53738_20514# a_54504_20259# 0.47248f
C915 a_53968_20434# a_53899_20488# 0.70262f
C916 a_58734_56203# VDD 0.35557f
C917 vco_wob_0.vctl m6_60810_42209# 0.05504f
C918 3bit_freq_divider_0.dff_nclk_0.nCLK a_53968_22190# 0.32534f
C919 a_53738_22270# VDD 0.21577f
C920 a_54434_21392# a_54472_21129# 0.36535f
C921 a_57173_40413# VDD 0.98193f
C922 a_55862_56737# charge_pump_0.bias_p 0.3307f
C923 3bit_freq_divider_1.dff_nclk_0.nCLK a_62900_21935# 0.27425f
C924 a_61887_24046# VDD 0.22153f
C925 3bit_freq_divider_1.dff_nclk_0.nCLK 3bit_freq_divider_1.freq_div_cell_0.Cout 0.32366f
C926 a_54504_22015# VDD 0.38024f
C927 a_53022_43738# a_55742_43159# 0.19603f
C928 a_53065_23691# VDD 0.44373f
C929 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.nQ 3bit_freq_divider_0.dff_nclk_0.nCLK 0.02505f
C930 a_61887_20534# a_62270_20543# 0.66077f
C931 a_61691_20534# a_62654_20215# 0.02302f
C932 a_59799_40285# VDD 1.38295f
C933 3bit_freq_divider_0.dff_nclk_0.D a_51693_23426# 0.04146f
C934 VDD Y2 1.18034f
C935 a_61707_25000# a_61675_24642# 0.0104f
C936 3bit_freq_divider_0.freq_div_cell_0.Cin 3bit_freq_divider_0.dff_nclk_0.nCLK 0.32366f
C937 a_53022_43738# a_57178_43159# 0.04298f
C938 a_60385_24717# a_60385_24558# 0.01952f
C939 vco_wob_0.vctl a_55969_42591# 0.0811f
C940 a_56039_25022# VDD 0.01215f
C941 a_54400_43159# a_54494_43159# 0.42202f
C942 m2_17285_2698# m3_17285_2698# 0.20496p
C943 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.Q X1 0.15458f
C944 a_51631_22774# a_51693_23075# 0.04255f
C945 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.Q a_61878_21130# 0.02559f
C946 a_60967_23234# VDD 0.45855f
C947 m1_17285_2698# CLK_IN 0.01061f
C948 3bit_freq_divider_0.dff_nclk_0.nRST X1 0.08188f
C949 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.D a_54504_23771# 0.3562f
C950 vco_wob_0.vctl a_58454_40850# 0.04998f
C951 a_54494_43159# a_55836_43159# 0.88103f
C952 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.Q 3bit_freq_divider_1.freq_div_cell_0.Cin 0.22232f
C953 charge_pump_0.vout a_54842_49733# 0.02265f
C954 a_62654_20215# 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.nQ 0.0571f
C955 3bit_freq_divider_1.dff_nclk_0.nCLK a_61394_20220# 0.37259f
C956 a_52886_24904# 3bit_freq_divider_0.sg13g2_or3_1_0.C 0.23357f
C957 a_51759_25014# a_51721_24988# 0.10864f
C958 PFD_0.VCO_CLK X0 0.1115f
C959 3bit_freq_divider_0.dff_nclk_0.nCLK a_53445_20214# 0.26292f
C960 3bit_freq_divider_1.freq_div_cell_1.Cout 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.D 0.04623f
C961 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.Q a_63255_23244# 0.12248f
C962 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.nQ Y1 0.01108f
C963 a_54434_24904# a_54472_24641# 0.36535f
C964 3bit_freq_divider_1.dff_nclk_0.nCLK a_63463_20216# 0.05882f
C965 PFD_0.UP CLK_IN 0.15472f
C966 a_54434_21392# 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.D 0.24715f
C967 3bit_freq_divider_1.sg13g2_or3_1_0.A Y2 0.10441f
C968 3bit_freq_divider_0.dff_nclk_0.D a_51684_22692# 0.0175f
C969 3bit_freq_divider_1.sg13g2_nand2_1_0.Y VDD 3.38844f
C970 3bit_freq_divider_0.dff_nclk_0.nCLK 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.60301f
C971 a_56013_24979# a_56038_24617# 0.01952f
C972 a_55742_43159# VDD 1.36686f
C973 a_62119_20605# VDD 0.2982f
C974 3bit_freq_divider_0.dff_nclk_0.nRST a_51684_22284# 0.34874f
C975 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 3bit_freq_divider_0.sg13g2_nand2_1_0.Y 0.1064f
C976 a_55345_23141# VDD 0.45855f
C977 a_57178_43159# VDD 1.11494f
C978 3bit_freq_divider_1.sg13g2_nand2_1_0.Y 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.11142f
C979 3bit_freq_divider_1.dff_nclk_0.nCLK 3bit_freq_divider_1.sg13g2_or3_1_0.B 0.58488f
C980 VDD X2 0.25402f
C981 3bit_freq_divider_1.sg13g2_tiehi_1.L_HI a_61707_25000# 0.12082f
C982 a_63255_25000# Y0 0.39999f
C983 a_64383_23628# a_64419_23326# 0.04304f
C984 a_52886_23148# a_52924_22885# 0.36535f
C985 a_60385_24947# VDD 0.11858f
C986 PFD_0.VCO_CLK a_51622_24863# 0.02673f
C987 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.Q Y1 0.15164f
C988 3bit_freq_divider_1.sg13g2_nand2_1_0.Y a_60967_21478# 0.08797f
C989 a_63255_23244# VDD 0.25835f
C990 m4_17285_2698# CLK_OUT 0.3817f
C991 a_48909_28913# CLK_IN 0.12375f
C992 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.D a_61691_24046# 0.01446f
C993 3bit_freq_divider_1.freq_div_cell_0.Cout 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.D 0.084f
C994 3bit_freq_divider_1.dff_nclk_0.nCLK 3bit_freq_divider_1.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.10701f
C995 a_51685_23725# VDD 0.30547f
C996 a_55345_21385# VDD 0.45855f
C997 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.sg13g2_dfrbp_1_0.CLK a_61887_24046# 0.01324f
C998 3bit_freq_divider_1.sg13g2_or3_1_0.C 3bit_freq_divider_1.sg13g2_or3_1_0.B 1.00414f
C999 a_53086_40850# a_53147_40413# 0.04971f
C1000 3bit_freq_divider_0.sg13g2_tiehi_1.L_HI a_56013_24979# 0.02161f
C1001 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.Q a_52924_24641# 0.02246f
C1002 a_54434_24904# 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.D 0.24715f
C1003 a_63255_23244# a_63223_22886# 0.0104f
C1004 charge_pump_0.bias_p a_56742_53480# 0.04781f
C1005 charge_pump_0.bias_n a_56828_53480# 0.01798f
C1006 a_56013_24979# a_55941_24882# 0.14868f
C1007 a_53147_40413# a_54489_40413# 0.35714f
C1008 a_58454_40850# a_57173_40413# 0.22936f
C1009 a_53738_22270# a_53968_22190# 0.13068f
C1010 3bit_freq_divider_0.EN VDD 6.40652f
C1011 3bit_freq_divider_1.dff_nclk_0.D a_64424_22200# 0.43097f
C1012 a_54472_22885# VDD 0.21321f
C1013 3bit_freq_divider_0.sg13g2_or3_1_0.C a_51693_23075# 0.01089f
C1014 a_61691_24046# a_61394_23732# 0.17766f
C1015 a_54489_40413# a_55769_40283# 0.45379f
C1016 a_55862_56737# a_55948_56737# 0.0609f
C1017 3bit_freq_divider_0.dff_nclk_0.nCLK 3bit_freq_divider_0.sg13g2_or3_1_0.B 0.58488f
C1018 a_53968_22190# a_54504_22015# 0.45825f
C1019 a_53774_20178# a_53899_20488# 0.04304f
C1020 VDD Y1 0.44908f
C1021 3bit_freq_divider_1.sg13g2_or3_1_0.C 3bit_freq_divider_1.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.28129f
C1022 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.Q a_61878_24642# 0.02559f
C1023 a_53065_21935# VDD 0.43552f
C1024 a_61887_24046# a_62119_24117# 0.13068f
C1025 a_64384_24445# a_64383_23889# 0.09575f
C1026 3bit_freq_divider_0.sg13g2_tiehi_1.L_HI a_54472_24641# 0.01011f
C1027 a_51759_25014# 3bit_freq_divider_0.dff_nclk_0.nRST 0.03098f
C1028 a_51721_24988# a_51622_24863# 0.0229f
C1029 a_54357_49278# VDD 0.31963f
C1030 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.D 3bit_freq_divider_0.sg13g2_nand2_1_0.Y 0.04726f
C1031 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.Q a_62654_20215# 0.01984f
C1032 a_64384_24445# CLK_OUT 0.1244f
C1033 a_54357_49278# PFD_0.DOWN 0.04759f
C1034 3bit_freq_divider_1.freq_div_cell_0.Cout a_61707_21488# 0.12082f
C1035 a_62654_23727# a_63463_23728# 0.09575f
C1036 3bit_freq_divider_1.dff_nclk_0.nRST a_64383_23300# 0.31482f
C1037 a_61887_22290# a_62270_22299# 0.66077f
C1038 m4_17285_2698# Y0 0.3817f
C1039 a_54472_21129# VDD 0.21321f
C1040 a_53065_23691# 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.nQ 0.05822f
C1041 a_61691_22290# a_62654_21971# 0.02302f
C1042 a_64383_23434# a_64383_23300# 0.13068f
C1043 a_51648_24438# VDD 0.24104f
C1044 3bit_freq_divider_1.sg13g2_nand2_1_0.Y 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.1064f
C1045 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.Q a_55345_24897# 0.30546f
C1046 a_57178_43159# m6_60810_42209# 0.08511f
C1047 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.Q 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.nQ 0.02712f
C1048 a_63463_23728# 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.nQ 0.21609f
C1049 a_53774_23690# a_53968_23946# 0.05314f
C1050 a_63463_21972# Y2 0.01788f
C1051 3bit_freq_divider_0.dff_nclk_0.nCLK 3bit_freq_divider_0.sg13g2_or3_1_0.A 0.48568f
C1052 a_52886_21392# VDD 0.26051f
C1053 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.D VDD 0.97883f
C1054 a_53022_43738# a_53086_40850# 0.06371f
C1055 a_53738_24026# a_53899_24000# 0.66077f
C1056 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.Q X2 0.17317f
C1057 a_62654_21971# 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.nQ 0.0571f
C1058 3bit_freq_divider_0.sg13g2_or3_1_0.C a_52924_24641# 0.10662f
C1059 a_56742_53480# nEN 0.28042f
C1060 3bit_freq_divider_1.sg13g2_or3_1_0.C 3bit_freq_divider_1.dff_nclk_0.nRST 0.57774f
C1061 3bit_freq_divider_1.sg13g2_or3_1_0.C a_64383_23434# 0.03556f
C1062 a_55836_43159# a_57311_42591# 0.03153f
C1063 a_53022_43738# a_54489_40413# 0.05403f
C1064 a_55941_24882# a_56137_24678# 0.0229f
C1065 a_51708_21299# VDD 0.01263f
C1066 3bit_freq_divider_0.sg13g2_or3_1_0.B 3bit_freq_divider_0.sg13g2_or3_1_0.A 0.72102f
C1067 a_53022_43738# a_57111_40283# 0.18962f
C1068 a_51685_23725# a_51684_22692# 0.04306f
C1069 VDD X1 1.47452f
C1070 3bit_freq_divider_0.dff_nclk_0.D 3bit_freq_divider_0.dff_nclk_0.nCLK 0.04354f
C1071 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.D VDD 0.9437f
C1072 3bit_freq_divider_1.freq_div_cell_0.Cin a_60967_23234# 0.13034f
C1073 3bit_freq_divider_0.CLK_IN a_58515_40413# 0.83094f
C1074 3bit_freq_divider_0.dff_nclk_0.nRST X0 0.14477f
C1075 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.Q a_55345_21385# 0.30546f
C1076 PFD_0.UP VDD 0.82664f
C1077 3bit_freq_divider_0.freq_div_cell_0.Cout 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.01369f
C1078 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.D a_61878_22886# 0.12185f
C1079 PFD_0.UP PFD_0.DOWN 0.20773f
C1080 m4_17285_2698# X0 0.39515f
C1081 m3_17285_2698# Y1 0.2919f
C1082 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.D VDD 0.97083f
R0 X1.n3 X1.n0 15.1893
R1 X1.n2 X1.n1 15.0005
R2 X1 X1.n3 9.55138
R3 X1.n1299 X1.n73 2.2505
R4 X1.n1303 X1.n70 2.2505
R5 X1.n1305 X1.n68 2.2505
R6 X1.n1309 X1.n65 2.2505
R7 X1.n1311 X1.n63 2.2505
R8 X1.n1315 X1.n60 2.2505
R9 X1.n1317 X1.n58 2.2505
R10 X1.n96 X1.n56 2.2505
R11 X1.n1322 X1.n54 2.2505
R12 X1.n158 X1.n51 2.2505
R13 X1.n1328 X1.n49 2.2505
R14 X1.n134 X1.n46 2.2505
R15 X1.n1334 X1.n44 2.2505
R16 X1.n112 X1.n40 2.2505
R17 X1.n37 X1.n28 2.2505
R18 X1.n1300 X1.n1299 2.2505
R19 X1.n1303 X1.n1302 2.2505
R20 X1.n1306 X1.n1305 2.2505
R21 X1.n1309 X1.n1308 2.2505
R22 X1.n1312 X1.n1311 2.2505
R23 X1.n1315 X1.n1314 2.2505
R24 X1.n1318 X1.n1317 2.2505
R25 X1.n1319 X1.n56 2.2505
R26 X1.n1322 X1.n52 2.2505
R27 X1.n1325 X1.n51 2.2505
R28 X1.n1328 X1.n47 2.2505
R29 X1.n1331 X1.n46 2.2505
R30 X1.n1334 X1.n42 2.2505
R31 X1.n1337 X1.n40 2.2505
R32 X1.n41 X1.n28 2.2505
R33 X1.n471 X1.n470 2.2505
R34 X1.n472 X1.n459 2.2505
R35 X1.n781 X1.n451 2.2505
R36 X1.n777 X1.n443 2.2505
R37 X1.n879 X1.n878 2.2505
R38 X1.n885 X1.n884 2.2505
R39 X1.n907 X1.n404 2.2505
R40 X1.n402 X1.n401 2.2505
R41 X1.n937 X1.n936 2.2505
R42 X1.n975 X1.n974 2.2505
R43 X1.n985 X1.n984 2.2505
R44 X1.n980 X1.n366 2.2505
R45 X1.n1026 X1.n351 2.2505
R46 X1.n1041 X1.n349 2.2505
R47 X1.n1073 X1.n337 2.2505
R48 X1.n775 X1.n471 2.2505
R49 X1.n784 X1.n472 2.2505
R50 X1.n781 X1.n776 2.2505
R51 X1.n778 X1.n777 2.2505
R52 X1.n880 X1.n879 2.2505
R53 X1.n884 X1.n883 2.2505
R54 X1.n404 X1.n403 2.2505
R55 X1.n934 X1.n402 2.2505
R56 X1.n936 X1.n935 2.2505
R57 X1.n976 X1.n975 2.2505
R58 X1.n984 X1.n983 2.2505
R59 X1.n981 X1.n980 2.2505
R60 X1.n351 X1.n350 2.2505
R61 X1.n1069 X1.n349 2.2505
R62 X1.n337 X1.n336 2.2505
R63 X1.n1286 X1.n74 2.2505
R64 X1.n1288 X1.n1287 2.2505
R65 X1.n1285 X1.n252 2.2505
R66 X1.n1284 X1.n1283 2.2505
R67 X1.n254 X1.n253 2.2505
R68 X1.n1263 X1.n1262 2.2505
R69 X1.n1261 X1.n261 2.2505
R70 X1.n1260 X1.n1259 2.2505
R71 X1.n263 X1.n262 2.2505
R72 X1.n1233 X1.n1232 2.2505
R73 X1.n1234 X1.n1231 2.2505
R74 X1.n1230 X1.n272 2.2505
R75 X1.n1229 X1.n1228 2.2505
R76 X1.n274 X1.n273 2.2505
R77 X1.n1209 X1.n1208 2.2505
R78 X1.n1207 X1.n282 2.2505
R79 X1.n1206 X1.n1205 2.2505
R80 X1.n284 X1.n283 2.2505
R81 X1.n1186 X1.n1185 2.2505
R82 X1.n1187 X1.n1184 2.2505
R83 X1.n1183 X1.n299 2.2505
R84 X1.n1182 X1.n1181 2.2505
R85 X1.n301 X1.n300 2.2505
R86 X1.n1155 X1.n1154 2.2505
R87 X1.n1156 X1.n1153 2.2505
R88 X1.n1152 X1.n311 2.2505
R89 X1.n1151 X1.n1150 2.2505
R90 X1.n313 X1.n312 2.2505
R91 X1.n1131 X1.n1130 2.2505
R92 X1.n1129 X1.n325 2.2505
R93 X1.n1128 X1.n1127 2.2505
R94 X1.n327 X1.n326 2.2505
R95 X1.n1109 X1.n1108 2.2505
R96 X1.n1107 X1.n335 2.2505
R97 X1.n1093 X1.n335 2.2505
R98 X1.n1110 X1.n1109 2.2505
R99 X1.n1113 X1.n327 2.2505
R100 X1.n1127 X1.n1126 2.2505
R101 X1.n329 X1.n325 2.2505
R102 X1.n1132 X1.n1131 2.2505
R103 X1.n1135 X1.n313 2.2505
R104 X1.n1150 X1.n1149 2.2505
R105 X1.n317 X1.n311 2.2505
R106 X1.n1157 X1.n1156 2.2505
R107 X1.n1155 X1.n308 2.2505
R108 X1.n1165 X1.n301 2.2505
R109 X1.n1181 X1.n1180 2.2505
R110 X1.n1170 X1.n299 2.2505
R111 X1.n1188 X1.n1187 2.2505
R112 X1.n1186 X1.n296 2.2505
R113 X1.n1196 X1.n284 2.2505
R114 X1.n1205 X1.n1204 2.2505
R115 X1.n290 X1.n282 2.2505
R116 X1.n1210 X1.n1209 2.2505
R117 X1.n1212 X1.n274 2.2505
R118 X1.n1228 X1.n1227 2.2505
R119 X1.n1217 X1.n272 2.2505
R120 X1.n1235 X1.n1234 2.2505
R121 X1.n1233 X1.n269 2.2505
R122 X1.n1243 X1.n263 2.2505
R123 X1.n1259 X1.n1258 2.2505
R124 X1.n1252 X1.n261 2.2505
R125 X1.n1264 X1.n1263 2.2505
R126 X1.n1267 X1.n254 2.2505
R127 X1.n1283 X1.n1282 2.2505
R128 X1.n1275 X1.n252 2.2505
R129 X1.n1289 X1.n1288 2.2505
R130 X1.n76 X1.n74 2.2505
R131 X1.n772 X1.n475 2.2505
R132 X1.n771 X1.n476 2.2505
R133 X1.n564 X1.n477 2.2505
R134 X1.n767 X1.n479 2.2505
R135 X1.n766 X1.n480 2.2505
R136 X1.n765 X1.n481 2.2505
R137 X1.n516 X1.n482 2.2505
R138 X1.n761 X1.n484 2.2505
R139 X1.n760 X1.n485 2.2505
R140 X1.n759 X1.n486 2.2505
R141 X1.n507 X1.n487 2.2505
R142 X1.n755 X1.n489 2.2505
R143 X1.n754 X1.n490 2.2505
R144 X1.n753 X1.n491 2.2505
R145 X1.n618 X1.n492 2.2505
R146 X1.n749 X1.n748 2.2505
R147 X1.n738 X1.n6 2.2505
R148 X1.n1374 X1.n7 2.2505
R149 X1.n1373 X1.n8 2.2505
R150 X1.n1372 X1.n9 2.2505
R151 X1.n630 X1.n10 2.2505
R152 X1.n1368 X1.n12 2.2505
R153 X1.n1367 X1.n13 2.2505
R154 X1.n1366 X1.n14 2.2505
R155 X1.n638 X1.n15 2.2505
R156 X1.n1362 X1.n17 2.2505
R157 X1.n1361 X1.n18 2.2505
R158 X1.n1360 X1.n19 2.2505
R159 X1.n689 X1.n20 2.2505
R160 X1.n1356 X1.n22 2.2505
R161 X1.n1355 X1.n23 2.2505
R162 X1.n1354 X1.n24 2.2505
R163 X1.n671 X1.n25 2.2505
R164 X1.n1350 X1.n27 2.2505
R165 X1.n1351 X1.n1350 2.2505
R166 X1.n1352 X1.n25 2.2505
R167 X1.n1354 X1.n1353 2.2505
R168 X1.n1355 X1.n21 2.2505
R169 X1.n1357 X1.n1356 2.2505
R170 X1.n1358 X1.n20 2.2505
R171 X1.n1360 X1.n1359 2.2505
R172 X1.n1361 X1.n16 2.2505
R173 X1.n1363 X1.n1362 2.2505
R174 X1.n1364 X1.n15 2.2505
R175 X1.n1366 X1.n1365 2.2505
R176 X1.n1367 X1.n11 2.2505
R177 X1.n1369 X1.n1368 2.2505
R178 X1.n1370 X1.n10 2.2505
R179 X1.n1372 X1.n1371 2.2505
R180 X1.n1373 X1.n5 2.2505
R181 X1.n1375 X1.n1374 2.2505
R182 X1.n6 X1.n4 2.2505
R183 X1.n750 X1.n749 2.2505
R184 X1.n751 X1.n492 2.2505
R185 X1.n753 X1.n752 2.2505
R186 X1.n754 X1.n488 2.2505
R187 X1.n756 X1.n755 2.2505
R188 X1.n757 X1.n487 2.2505
R189 X1.n759 X1.n758 2.2505
R190 X1.n760 X1.n483 2.2505
R191 X1.n762 X1.n761 2.2505
R192 X1.n763 X1.n482 2.2505
R193 X1.n765 X1.n764 2.2505
R194 X1.n766 X1.n478 2.2505
R195 X1.n768 X1.n767 2.2505
R196 X1.n769 X1.n477 2.2505
R197 X1.n771 X1.n770 2.2505
R198 X1.n772 X1.n473 2.2505
R199 X1.n77 X1.n75 2.2005
R200 X1.n34 X1.n29 2.2005
R201 X1.n38 X1.n35 2.2005
R202 X1.n1342 X1.n1341 2.2005
R203 X1.n39 X1.n36 2.2005
R204 X1.n115 X1.n114 2.2005
R205 X1.n117 X1.n116 2.2005
R206 X1.n119 X1.n118 2.2005
R207 X1.n121 X1.n120 2.2005
R208 X1.n123 X1.n122 2.2005
R209 X1.n125 X1.n124 2.2005
R210 X1.n127 X1.n126 2.2005
R211 X1.n129 X1.n128 2.2005
R212 X1.n132 X1.n131 2.2005
R213 X1.n133 X1.n107 2.2005
R214 X1.n137 X1.n136 2.2005
R215 X1.n135 X1.n105 2.2005
R216 X1.n143 X1.n142 2.2005
R217 X1.n144 X1.n104 2.2005
R218 X1.n146 X1.n145 2.2005
R219 X1.n149 X1.n148 2.2005
R220 X1.n151 X1.n150 2.2005
R221 X1.n102 X1.n101 2.2005
R222 X1.n157 X1.n156 2.2005
R223 X1.n159 X1.n100 2.2005
R224 X1.n161 X1.n160 2.2005
R225 X1.n163 X1.n162 2.2005
R226 X1.n165 X1.n164 2.2005
R227 X1.n167 X1.n166 2.2005
R228 X1.n170 X1.n169 2.2005
R229 X1.n168 X1.n97 2.2005
R230 X1.n177 X1.n176 2.2005
R231 X1.n179 X1.n178 2.2005
R232 X1.n181 X1.n180 2.2005
R233 X1.n183 X1.n182 2.2005
R234 X1.n185 X1.n184 2.2005
R235 X1.n187 X1.n186 2.2005
R236 X1.n189 X1.n188 2.2005
R237 X1.n191 X1.n190 2.2005
R238 X1.n194 X1.n193 2.2005
R239 X1.n195 X1.n93 2.2005
R240 X1.n199 X1.n198 2.2005
R241 X1.n197 X1.n91 2.2005
R242 X1.n205 X1.n204 2.2005
R243 X1.n206 X1.n90 2.2005
R244 X1.n208 X1.n207 2.2005
R245 X1.n211 X1.n210 2.2005
R246 X1.n213 X1.n212 2.2005
R247 X1.n88 X1.n87 2.2005
R248 X1.n221 X1.n220 2.2005
R249 X1.n223 X1.n86 2.2005
R250 X1.n225 X1.n224 2.2005
R251 X1.n227 X1.n226 2.2005
R252 X1.n229 X1.n228 2.2005
R253 X1.n231 X1.n230 2.2005
R254 X1.n233 X1.n232 2.2005
R255 X1.n235 X1.n234 2.2005
R256 X1.n237 X1.n83 2.2005
R257 X1.n239 X1.n238 2.2005
R258 X1.n241 X1.n82 2.2005
R259 X1.n243 X1.n242 2.2005
R260 X1.n1083 X1.n338 2.2005
R261 X1.n1074 X1.n345 2.2005
R262 X1.n1076 X1.n1075 2.2005
R263 X1.n1048 X1.n348 2.2005
R264 X1.n1053 X1.n1043 2.2005
R265 X1.n1042 X1.n1039 2.2005
R266 X1.n1060 X1.n353 2.2005
R267 X1.n1065 X1.n1064 2.2005
R268 X1.n1035 X1.n352 2.2005
R269 X1.n1033 X1.n358 2.2005
R270 X1.n1028 X1.n1027 2.2005
R271 X1.n1025 X1.n1024 2.2005
R272 X1.n1018 X1.n1017 2.2005
R273 X1.n1016 X1.n1015 2.2005
R274 X1.n1010 X1.n1009 2.2005
R275 X1.n1008 X1.n1007 2.2005
R276 X1.n1002 X1.n1001 2.2005
R277 X1.n1000 X1.n999 2.2005
R278 X1.n993 X1.n375 2.2005
R279 X1.n987 X1.n986 2.2005
R280 X1.n381 X1.n380 2.2005
R281 X1.n967 X1.n388 2.2005
R282 X1.n973 X1.n972 2.2005
R283 X1.n961 X1.n386 2.2005
R284 X1.n955 X1.n954 2.2005
R285 X1.n952 X1.n951 2.2005
R286 X1.n947 X1.n395 2.2005
R287 X1.n938 X1.n398 2.2005
R288 X1.n940 X1.n939 2.2005
R289 X1.n924 X1.n406 2.2005
R290 X1.n930 X1.n929 2.2005
R291 X1.n917 X1.n405 2.2005
R292 X1.n908 X1.n410 2.2005
R293 X1.n910 X1.n909 2.2005
R294 X1.n906 X1.n905 2.2005
R295 X1.n899 X1.n413 2.2005
R296 X1.n425 X1.n417 2.2005
R297 X1.n892 X1.n420 2.2005
R298 X1.n887 X1.n886 2.2005
R299 X1.n870 X1.n423 2.2005
R300 X1.n434 X1.n432 2.2005
R301 X1.n877 X1.n876 2.2005
R302 X1.n863 X1.n430 2.2005
R303 X1.n857 X1.n856 2.2005
R304 X1.n855 X1.n854 2.2005
R305 X1.n849 X1.n848 2.2005
R306 X1.n847 X1.n846 2.2005
R307 X1.n842 X1.n841 2.2005
R308 X1.n840 X1.n839 2.2005
R309 X1.n833 X1.n832 2.2005
R310 X1.n831 X1.n830 2.2005
R311 X1.n823 X1.n822 2.2005
R312 X1.n821 X1.n820 2.2005
R313 X1.n814 X1.n813 2.2005
R314 X1.n812 X1.n811 2.2005
R315 X1.n806 X1.n805 2.2005
R316 X1.n804 X1.n803 2.2005
R317 X1.n797 X1.n463 2.2005
R318 X1.n788 X1.n467 2.2005
R319 X1.n790 X1.n789 2.2005
R320 X1.n538 X1.n536 2.2005
R321 X1.n1091 X1.n339 2.2005
R322 X1.n1095 X1.n1094 2.2005
R323 X1.n1096 X1.n334 2.2005
R324 X1.n1111 X1.n332 2.2005
R325 X1.n1115 X1.n1114 2.2005
R326 X1.n1112 X1.n333 2.2005
R327 X1.n330 X1.n328 2.2005
R328 X1.n1125 X1.n1124 2.2005
R329 X1.n1123 X1.n1122 2.2005
R330 X1.n1120 X1.n324 2.2005
R331 X1.n1133 X1.n321 2.2005
R332 X1.n1137 X1.n1136 2.2005
R333 X1.n1134 X1.n323 2.2005
R334 X1.n322 X1.n314 2.2005
R335 X1.n1148 X1.n1147 2.2005
R336 X1.n1146 X1.n315 2.2005
R337 X1.n319 X1.n318 2.2005
R338 X1.n1141 X1.n310 2.2005
R339 X1.n1158 X1.n309 2.2005
R340 X1.n1160 X1.n1159 2.2005
R341 X1.n1163 X1.n1162 2.2005
R342 X1.n1164 X1.n307 2.2005
R343 X1.n1167 X1.n1166 2.2005
R344 X1.n304 X1.n302 2.2005
R345 X1.n1179 X1.n1178 2.2005
R346 X1.n305 X1.n303 2.2005
R347 X1.n1172 X1.n1171 2.2005
R348 X1.n1173 X1.n298 2.2005
R349 X1.n1189 X1.n297 2.2005
R350 X1.n1191 X1.n1190 2.2005
R351 X1.n1194 X1.n1193 2.2005
R352 X1.n1195 X1.n295 2.2005
R353 X1.n1198 X1.n1197 2.2005
R354 X1.n287 X1.n285 2.2005
R355 X1.n1203 X1.n1202 2.2005
R356 X1.n293 X1.n286 2.2005
R357 X1.n292 X1.n291 2.2005
R358 X1.n288 X1.n281 2.2005
R359 X1.n1211 X1.n280 2.2005
R360 X1.n1214 X1.n1213 2.2005
R361 X1.n277 X1.n275 2.2005
R362 X1.n1226 X1.n1225 2.2005
R363 X1.n278 X1.n276 2.2005
R364 X1.n1219 X1.n1218 2.2005
R365 X1.n1220 X1.n271 2.2005
R366 X1.n1236 X1.n270 2.2005
R367 X1.n1238 X1.n1237 2.2005
R368 X1.n1241 X1.n1240 2.2005
R369 X1.n1242 X1.n268 2.2005
R370 X1.n1245 X1.n1244 2.2005
R371 X1.n266 X1.n264 2.2005
R372 X1.n1257 X1.n1256 2.2005
R373 X1.n1255 X1.n265 2.2005
R374 X1.n1254 X1.n1253 2.2005
R375 X1.n1250 X1.n260 2.2005
R376 X1.n1265 X1.n259 2.2005
R377 X1.n1269 X1.n1268 2.2005
R378 X1.n1266 X1.n257 2.2005
R379 X1.n1274 X1.n255 2.2005
R380 X1.n1281 X1.n1280 2.2005
R381 X1.n1279 X1.n256 2.2005
R382 X1.n1277 X1.n1276 2.2005
R383 X1.n251 X1.n250 2.2005
R384 X1.n1292 X1.n1291 2.2005
R385 X1.n1290 X1.n78 2.2005
R386 X1.n549 X1.n548 2.2005
R387 X1.n553 X1.n552 2.2005
R388 X1.n551 X1.n526 2.2005
R389 X1.n560 X1.n558 2.2005
R390 X1.n566 X1.n565 2.2005
R391 X1.n563 X1.n559 2.2005
R392 X1.n562 X1.n561 2.2005
R393 X1.n523 X1.n522 2.2005
R394 X1.n575 X1.n570 2.2005
R395 X1.n577 X1.n576 2.2005
R396 X1.n573 X1.n572 2.2005
R397 X1.n571 X1.n517 2.2005
R398 X1.n584 X1.n583 2.2005
R399 X1.n586 X1.n585 2.2005
R400 X1.n589 X1.n588 2.2005
R401 X1.n591 X1.n590 2.2005
R402 X1.n595 X1.n594 2.2005
R403 X1.n593 X1.n592 2.2005
R404 X1.n512 X1.n511 2.2005
R405 X1.n510 X1.n508 2.2005
R406 X1.n603 X1.n602 2.2005
R407 X1.n605 X1.n604 2.2005
R408 X1.n607 X1.n606 2.2005
R409 X1.n609 X1.n608 2.2005
R410 X1.n611 X1.n610 2.2005
R411 X1.n613 X1.n612 2.2005
R412 X1.n616 X1.n615 2.2005
R413 X1.n617 X1.n501 2.2005
R414 X1.n620 X1.n619 2.2005
R415 X1.n502 X1.n493 2.2005
R416 X1.n747 X1.n746 2.2005
R417 X1.n745 X1.n494 2.2005
R418 X1.n739 X1.n496 2.2005
R419 X1.n741 X1.n740 2.2005
R420 X1.n736 X1.n735 2.2005
R421 X1.n734 X1.n733 2.2005
R422 X1.n731 X1.n730 2.2005
R423 X1.n729 X1.n728 2.2005
R424 X1.n727 X1.n726 2.2005
R425 X1.n725 X1.n724 2.2005
R426 X1.n722 X1.n721 2.2005
R427 X1.n714 X1.n633 2.2005
R428 X1.n716 X1.n715 2.2005
R429 X1.n712 X1.n711 2.2005
R430 X1.n710 X1.n709 2.2005
R431 X1.n707 X1.n706 2.2005
R432 X1.n705 X1.n704 2.2005
R433 X1.n702 X1.n701 2.2005
R434 X1.n700 X1.n699 2.2005
R435 X1.n641 X1.n640 2.2005
R436 X1.n643 X1.n642 2.2005
R437 X1.n647 X1.n646 2.2005
R438 X1.n649 X1.n648 2.2005
R439 X1.n686 X1.n685 2.2005
R440 X1.n688 X1.n687 2.2005
R441 X1.n690 X1.n653 2.2005
R442 X1.n692 X1.n691 2.2005
R443 X1.n684 X1.n683 2.2005
R444 X1.n682 X1.n681 2.2005
R445 X1.n660 X1.n658 2.2005
R446 X1.n662 X1.n661 2.2005
R447 X1.n674 X1.n673 2.2005
R448 X1.n672 X1.n664 2.2005
R449 X1.n670 X1.n669 2.2005
R450 X1.n668 X1.n665 2.2005
R451 X1.n240 X1.n71 1.8005
R452 X1.n1304 X1.n69 1.8005
R453 X1.n222 X1.n66 1.8005
R454 X1.n1310 X1.n64 1.8005
R455 X1.n196 X1.n61 1.8005
R456 X1.n1316 X1.n59 1.8005
R457 X1.n1321 X1.n55 1.8005
R458 X1.n1323 X1.n53 1.8005
R459 X1.n1327 X1.n50 1.8005
R460 X1.n1329 X1.n48 1.8005
R461 X1.n1333 X1.n45 1.8005
R462 X1.n1335 X1.n43 1.8005
R463 X1.n1340 X1.n1339 1.8005
R464 X1.n1301 X1.n71 1.8005
R465 X1.n1304 X1.n67 1.8005
R466 X1.n1307 X1.n66 1.8005
R467 X1.n1310 X1.n62 1.8005
R468 X1.n1313 X1.n61 1.8005
R469 X1.n1316 X1.n57 1.8005
R470 X1.n1321 X1.n1320 1.8005
R471 X1.n1324 X1.n1323 1.8005
R472 X1.n1327 X1.n1326 1.8005
R473 X1.n1330 X1.n1329 1.8005
R474 X1.n1333 X1.n1332 1.8005
R475 X1.n1336 X1.n1335 1.8005
R476 X1.n1339 X1.n1338 1.8005
R477 X1.n787 X1.n786 1.8005
R478 X1.n782 X1.n455 1.8005
R479 X1.n780 X1.n447 1.8005
R480 X1.n439 X1.n429 1.8005
R481 X1.n431 X1.n424 1.8005
R482 X1.n427 X1.n426 1.8005
R483 X1.n932 X1.n931 1.8005
R484 X1.n953 X1.n385 1.8005
R485 X1.n387 X1.n382 1.8005
R486 X1.n383 X1.n371 1.8005
R487 X1.n979 X1.n361 1.8005
R488 X1.n1067 X1.n1066 1.8005
R489 X1.n1072 X1.n1071 1.8005
R490 X1.n786 X1.n785 1.8005
R491 X1.n783 X1.n782 1.8005
R492 X1.n780 X1.n779 1.8005
R493 X1.n429 X1.n428 1.8005
R494 X1.n881 X1.n424 1.8005
R495 X1.n882 X1.n427 1.8005
R496 X1.n933 X1.n932 1.8005
R497 X1.n385 X1.n384 1.8005
R498 X1.n977 X1.n382 1.8005
R499 X1.n982 X1.n383 1.8005
R500 X1.n979 X1.n978 1.8005
R501 X1.n1068 X1.n1067 1.8005
R502 X1.n1071 X1.n1070 1.8005
R503 X1.n1298 X1.n72 1.8005
R504 X1.n1298 X1.n1297 1.8005
R505 X1.n1349 X1.n1348 1.8005
R506 X1.n1349 X1.n26 1.8005
R507 X1.n1106 X1.n1105 1.5005
R508 X1.n1105 X1.n1104 1.5005
R509 X1.n773 X1.n474 1.5005
R510 X1.n774 X1.n773 1.5005
R511 X1.n1100 X1.n1092 1.1125
R512 X1.n678 X1.n659 1.10836
R513 X1.n680 X1.n679 1.10443
R514 X1.n32 X1.n31 1.10381
R515 X1.n1101 X1.n342 1.10372
R516 X1.n654 X1.n652 1.10339
R517 X1.n674 X1.n663 1.10272
R518 X1.n677 X1.n662 1.10272
R519 X1.n681 X1.n657 1.10272
R520 X1.n1099 X1.n1095 1.10263
R521 X1.n1096 X1.n331 1.10263
R522 X1.n245 X1.n244 1.1005
R523 X1.n1344 X1.n1343 1.1005
R524 X1.n113 X1.n33 1.1005
R525 X1.n111 X1.n110 1.1005
R526 X1.n109 X1.n108 1.1005
R527 X1.n130 X1.n106 1.1005
R528 X1.n139 X1.n138 1.1005
R529 X1.n141 X1.n140 1.1005
R530 X1.n147 X1.n103 1.1005
R531 X1.n153 X1.n152 1.1005
R532 X1.n155 X1.n154 1.1005
R533 X1.n99 X1.n98 1.1005
R534 X1.n172 X1.n171 1.1005
R535 X1.n176 X1.n175 1.1005
R536 X1.n174 X1.n95 1.1005
R537 X1.n173 X1.n94 1.1005
R538 X1.n192 X1.n92 1.1005
R539 X1.n201 X1.n200 1.1005
R540 X1.n203 X1.n202 1.1005
R541 X1.n209 X1.n89 1.1005
R542 X1.n215 X1.n214 1.1005
R543 X1.n219 X1.n218 1.1005
R544 X1.n217 X1.n85 1.1005
R545 X1.n216 X1.n84 1.1005
R546 X1.n236 X1.n81 1.1005
R547 X1.n1345 X1.n30 1.1005
R548 X1.n80 X1.n79 1.1005
R549 X1.n248 X1.n247 1.1005
R550 X1.n247 X1.n246 1.1005
R551 X1.n1296 X1.n1295 1.1005
R552 X1.n1294 X1.n1293 1.1005
R553 X1.n1278 X1.n249 1.1005
R554 X1.n1273 X1.n1272 1.1005
R555 X1.n1271 X1.n1270 1.1005
R556 X1.n1251 X1.n258 1.1005
R557 X1.n1249 X1.n1248 1.1005
R558 X1.n1247 X1.n1246 1.1005
R559 X1.n1239 X1.n267 1.1005
R560 X1.n1222 X1.n1221 1.1005
R561 X1.n1224 X1.n1223 1.1005
R562 X1.n1216 X1.n1215 1.1005
R563 X1.n289 X1.n279 1.1005
R564 X1.n1201 X1.n1200 1.1005
R565 X1.n1199 X1.n1198 1.1005
R566 X1.n1192 X1.n294 1.1005
R567 X1.n1175 X1.n1174 1.1005
R568 X1.n1177 X1.n1176 1.1005
R569 X1.n1169 X1.n1168 1.1005
R570 X1.n1161 X1.n306 1.1005
R571 X1.n1143 X1.n1142 1.1005
R572 X1.n1145 X1.n1144 1.1005
R573 X1.n1140 X1.n316 1.1005
R574 X1.n1139 X1.n1138 1.1005
R575 X1.n1121 X1.n320 1.1005
R576 X1.n1119 X1.n1118 1.1005
R577 X1.n1117 X1.n1116 1.1005
R578 X1.n1098 X1.n1097 1.1005
R579 X1.n1090 X1.n341 1.1005
R580 X1.n1103 X1.n1102 1.1005
R581 X1.n1089 X1.n1088 1.1005
R582 X1.n1086 X1.n341 1.1005
R583 X1.n1084 X1.n1083 1.1005
R584 X1.n1081 X1.n1080 1.1005
R585 X1.n1079 X1.n345 1.1005
R586 X1.n1076 X1.n346 1.1005
R587 X1.n1047 X1.n1046 1.1005
R588 X1.n1051 X1.n1044 1.1005
R589 X1.n1053 X1.n1052 1.1005
R590 X1.n1054 X1.n1040 1.1005
R591 X1.n1059 X1.n1038 1.1005
R592 X1.n1034 X1.n356 1.1005
R593 X1.n1033 X1.n1032 1.1005
R594 X1.n1031 X1.n357 1.1005
R595 X1.n1022 X1.n363 1.1005
R596 X1.n1024 X1.n1023 1.1005
R597 X1.n1021 X1.n362 1.1005
R598 X1.n1013 X1.n368 1.1005
R599 X1.n1004 X1.n372 1.1005
R600 X1.n1003 X1.n1002 1.1005
R601 X1.n374 X1.n373 1.1005
R602 X1.n995 X1.n994 1.1005
R603 X1.n993 X1.n377 1.1005
R604 X1.n992 X1.n991 1.1005
R605 X1.n989 X1.n988 1.1005
R606 X1.n380 X1.n379 1.1005
R607 X1.n968 X1.n967 1.1005
R608 X1.n971 X1.n970 1.1005
R609 X1.n963 X1.n962 1.1005
R610 X1.n961 X1.n391 1.1005
R611 X1.n960 X1.n959 1.1005
R612 X1.n394 X1.n393 1.1005
R613 X1.n945 X1.n944 1.1005
R614 X1.n943 X1.n398 1.1005
R615 X1.n940 X1.n399 1.1005
R616 X1.n923 X1.n922 1.1005
R617 X1.n927 X1.n408 1.1005
R618 X1.n929 X1.n928 1.1005
R619 X1.n920 X1.n407 1.1005
R620 X1.n915 X1.n914 1.1005
R621 X1.n903 X1.n415 1.1005
R622 X1.n905 X1.n904 1.1005
R623 X1.n900 X1.n899 1.1005
R624 X1.n897 X1.n896 1.1005
R625 X1.n893 X1.n418 1.1005
R626 X1.n892 X1.n891 1.1005
R627 X1.n890 X1.n419 1.1005
R628 X1.n869 X1.n868 1.1005
R629 X1.n865 X1.n864 1.1005
R630 X1.n863 X1.n435 1.1005
R631 X1.n862 X1.n861 1.1005
R632 X1.n438 X1.n437 1.1005
R633 X1.n854 X1.n853 1.1005
R634 X1.n852 X1.n440 1.1005
R635 X1.n442 X1.n441 1.1005
R636 X1.n846 X1.n845 1.1005
R637 X1.n843 X1.n842 1.1005
R638 X1.n838 X1.n837 1.1005
R639 X1.n835 X1.n834 1.1005
R640 X1.n833 X1.n449 1.1005
R641 X1.n827 X1.n450 1.1005
R642 X1.n825 X1.n824 1.1005
R643 X1.n823 X1.n453 1.1005
R644 X1.n817 X1.n454 1.1005
R645 X1.n816 X1.n456 1.1005
R646 X1.n815 X1.n814 1.1005
R647 X1.n811 X1.n810 1.1005
R648 X1.n808 X1.n807 1.1005
R649 X1.n801 X1.n465 1.1005
R650 X1.n803 X1.n802 1.1005
R651 X1.n800 X1.n464 1.1005
R652 X1.n795 X1.n794 1.1005
R653 X1.n537 X1.n535 1.1005
R654 X1.n539 X1.n538 1.1005
R655 X1.n540 X1.n529 1.1005
R656 X1.n793 X1.n467 1.1005
R657 X1.n792 X1.n791 1.1005
R658 X1.n790 X1.n468 1.1005
R659 X1.n534 X1.n469 1.1005
R660 X1.n796 X1.n466 1.1005
R661 X1.n799 X1.n798 1.1005
R662 X1.n462 X1.n461 1.1005
R663 X1.n809 X1.n460 1.1005
R664 X1.n458 X1.n457 1.1005
R665 X1.n819 X1.n818 1.1005
R666 X1.n826 X1.n452 1.1005
R667 X1.n829 X1.n828 1.1005
R668 X1.n836 X1.n448 1.1005
R669 X1.n446 X1.n445 1.1005
R670 X1.n844 X1.n444 1.1005
R671 X1.n851 X1.n850 1.1005
R672 X1.n859 X1.n858 1.1005
R673 X1.n860 X1.n436 1.1005
R674 X1.n866 X1.n433 1.1005
R675 X1.n870 X1.n867 1.1005
R676 X1.n872 X1.n871 1.1005
R677 X1.n873 X1.n434 1.1005
R678 X1.n875 X1.n874 1.1005
R679 X1.n422 X1.n421 1.1005
R680 X1.n889 X1.n888 1.1005
R681 X1.n895 X1.n894 1.1005
R682 X1.n898 X1.n416 1.1005
R683 X1.n901 X1.n414 1.1005
R684 X1.n913 X1.n410 1.1005
R685 X1.n912 X1.n911 1.1005
R686 X1.n910 X1.n411 1.1005
R687 X1.n902 X1.n412 1.1005
R688 X1.n916 X1.n409 1.1005
R689 X1.n919 X1.n918 1.1005
R690 X1.n926 X1.n925 1.1005
R691 X1.n921 X1.n400 1.1005
R692 X1.n942 X1.n941 1.1005
R693 X1.n951 X1.n950 1.1005
R694 X1.n949 X1.n396 1.1005
R695 X1.n948 X1.n947 1.1005
R696 X1.n946 X1.n397 1.1005
R697 X1.n957 X1.n956 1.1005
R698 X1.n958 X1.n392 1.1005
R699 X1.n964 X1.n389 1.1005
R700 X1.n969 X1.n390 1.1005
R701 X1.n966 X1.n965 1.1005
R702 X1.n990 X1.n378 1.1005
R703 X1.n996 X1.n376 1.1005
R704 X1.n998 X1.n997 1.1005
R705 X1.n1006 X1.n1005 1.1005
R706 X1.n1015 X1.n1014 1.1005
R707 X1.n1012 X1.n367 1.1005
R708 X1.n1011 X1.n1010 1.1005
R709 X1.n370 X1.n369 1.1005
R710 X1.n365 X1.n364 1.1005
R711 X1.n1020 X1.n1019 1.1005
R712 X1.n360 X1.n359 1.1005
R713 X1.n1030 X1.n1029 1.1005
R714 X1.n1036 X1.n1035 1.1005
R715 X1.n1061 X1.n1060 1.1005
R716 X1.n1062 X1.n355 1.1005
R717 X1.n1064 X1.n1063 1.1005
R718 X1.n1037 X1.n354 1.1005
R719 X1.n1058 X1.n1057 1.1005
R720 X1.n1056 X1.n1055 1.1005
R721 X1.n1050 X1.n1049 1.1005
R722 X1.n1045 X1.n347 1.1005
R723 X1.n1078 X1.n1077 1.1005
R724 X1.n1088 X1.n1087 1.1005
R725 X1.n1082 X1.n344 1.1005
R726 X1.n1085 X1.n340 1.1005
R727 X1.n545 X1.n527 1.1005
R728 X1.n556 X1.n555 1.1005
R729 X1.n578 X1.n520 1.1005
R730 X1.n621 X1.n499 1.1005
R731 X1.n627 X1.n626 1.1005
R732 X1.n717 X1.n634 1.1005
R733 X1.n533 X1.n530 1.1005
R734 X1.n542 X1.n528 1.1005
R735 X1.n547 X1.n546 1.1005
R736 X1.n667 X1.n666 1.1005
R737 X1.n676 X1.n675 1.1005
R738 X1.n656 X1.n655 1.1005
R739 X1.n694 X1.n693 1.1005
R740 X1.n698 X1.n697 1.1005
R741 X1.n719 X1.n718 1.1005
R742 X1.n631 X1.n628 1.1005
R743 X1.n625 X1.n497 1.1005
R744 X1.n624 X1.n495 1.1005
R745 X1.n623 X1.n622 1.1005
R746 X1.n599 X1.n505 1.1005
R747 X1.n597 X1.n596 1.1005
R748 X1.n580 X1.n579 1.1005
R749 X1.n568 X1.n567 1.1005
R750 X1.n554 X1.n525 1.1005
R751 X1.n544 X1.n543 1.1005
R752 X1.n531 X1.n530 1.1005
R753 X1.n542 X1.n541 1.1005
R754 X1.n1297 X1.n1296 0.733833
R755 X1.n1104 X1.n1103 0.733833
R756 X1.n543 X1.n474 0.733833
R757 X1.n1348 X1.n1347 0.733833
R758 X1.n713 X1.n634 0.573769
R759 X1.n574 X1.n520 0.573769
R760 X1.n732 X1.n627 0.573695
R761 X1.n557 X1.n556 0.573695
R762 X1.n503 X1.n499 0.573346
R763 X1.n743 X1.n742 0.573297
R764 X1.n343 X1.n341 0.550549
R765 X1.n542 X1.n532 0.550549
R766 X1.n720 X1.n719 0.39244
R767 X1.n580 X1.n519 0.39244
R768 X1.n737 X1.n497 0.389994
R769 X1.n550 X1.n525 0.389994
R770 X1.n623 X1.n498 0.387191
R771 X1.n695 X1.n650 0.384705
R772 X1.n601 X1.n600 0.384705
R773 X1.n708 X1.n635 0.384705
R774 X1.n582 X1.n581 0.384705
R775 X1.n696 X1.n645 0.382331
R776 X1.n598 X1.n513 0.382331
R777 X1.n639 X1.n637 0.382034
R778 X1.n515 X1.n514 0.382034
R779 X1.n632 X1.n629 0.379547
R780 X1.n614 X1.n500 0.379547
R781 X1.n569 X1.n521 0.379547
R782 X1.n723 X1.n632 0.375976
R783 X1.n569 X1.n524 0.375976
R784 X1.n504 X1.n500 0.375884
R785 X1.n703 X1.n639 0.374982
R786 X1.n587 X1.n514 0.374982
R787 X1.n696 X1.n644 0.374889
R788 X1.n598 X1.n509 0.374889
R789 X1.n695 X1.n651 0.373984
R790 X1.n600 X1.n506 0.373984
R791 X1.n636 X1.n635 0.373891
R792 X1.n581 X1.n518 0.373891
R793 X1.n744 X1.n743 0.280767
R794 X1.n1347 X1.n1346 0.275034
R795 X1.n3 X1.n2 0.182739
R796 X1 X1.n1376 0.0685591
R797 X1.n2 X1 0.0563209
R798 X1.n1339 X1.n28 0.0405
R799 X1.n1339 X1.n40 0.0405
R800 X1.n1335 X1.n40 0.0405
R801 X1.n1335 X1.n1334 0.0405
R802 X1.n1334 X1.n1333 0.0405
R803 X1.n1333 X1.n46 0.0405
R804 X1.n1329 X1.n46 0.0405
R805 X1.n1329 X1.n1328 0.0405
R806 X1.n1328 X1.n1327 0.0405
R807 X1.n1327 X1.n51 0.0405
R808 X1.n1323 X1.n51 0.0405
R809 X1.n1323 X1.n1322 0.0405
R810 X1.n1322 X1.n1321 0.0405
R811 X1.n1321 X1.n56 0.0405
R812 X1.n1317 X1.n1316 0.0405
R813 X1.n1316 X1.n1315 0.0405
R814 X1.n1315 X1.n61 0.0405
R815 X1.n1311 X1.n61 0.0405
R816 X1.n1311 X1.n1310 0.0405
R817 X1.n1310 X1.n1309 0.0405
R818 X1.n1309 X1.n66 0.0405
R819 X1.n1305 X1.n66 0.0405
R820 X1.n1305 X1.n1304 0.0405
R821 X1.n1304 X1.n1303 0.0405
R822 X1.n1303 X1.n71 0.0405
R823 X1.n1299 X1.n71 0.0405
R824 X1.n1338 X1.n41 0.0405
R825 X1.n1338 X1.n1337 0.0405
R826 X1.n1337 X1.n1336 0.0405
R827 X1.n1336 X1.n42 0.0405
R828 X1.n1332 X1.n42 0.0405
R829 X1.n1332 X1.n1331 0.0405
R830 X1.n1331 X1.n1330 0.0405
R831 X1.n1330 X1.n47 0.0405
R832 X1.n1326 X1.n47 0.0405
R833 X1.n1326 X1.n1325 0.0405
R834 X1.n1325 X1.n1324 0.0405
R835 X1.n1324 X1.n52 0.0405
R836 X1.n1320 X1.n52 0.0405
R837 X1.n1320 X1.n1319 0.0405
R838 X1.n1318 X1.n57 0.0405
R839 X1.n1314 X1.n57 0.0405
R840 X1.n1314 X1.n1313 0.0405
R841 X1.n1313 X1.n1312 0.0405
R842 X1.n1312 X1.n62 0.0405
R843 X1.n1308 X1.n62 0.0405
R844 X1.n1308 X1.n1307 0.0405
R845 X1.n1307 X1.n1306 0.0405
R846 X1.n1306 X1.n67 0.0405
R847 X1.n1302 X1.n67 0.0405
R848 X1.n1302 X1.n1301 0.0405
R849 X1.n1301 X1.n1300 0.0405
R850 X1.n786 X1.n471 0.0405
R851 X1.n786 X1.n472 0.0405
R852 X1.n782 X1.n472 0.0405
R853 X1.n782 X1.n781 0.0405
R854 X1.n781 X1.n780 0.0405
R855 X1.n780 X1.n777 0.0405
R856 X1.n777 X1.n429 0.0405
R857 X1.n879 X1.n429 0.0405
R858 X1.n879 X1.n424 0.0405
R859 X1.n884 X1.n424 0.0405
R860 X1.n884 X1.n427 0.0405
R861 X1.n427 X1.n404 0.0405
R862 X1.n932 X1.n404 0.0405
R863 X1.n932 X1.n402 0.0405
R864 X1.n936 X1.n385 0.0405
R865 X1.n975 X1.n385 0.0405
R866 X1.n975 X1.n382 0.0405
R867 X1.n984 X1.n382 0.0405
R868 X1.n984 X1.n383 0.0405
R869 X1.n980 X1.n383 0.0405
R870 X1.n980 X1.n979 0.0405
R871 X1.n979 X1.n351 0.0405
R872 X1.n1067 X1.n351 0.0405
R873 X1.n1067 X1.n349 0.0405
R874 X1.n1071 X1.n349 0.0405
R875 X1.n1071 X1.n337 0.0405
R876 X1.n785 X1.n775 0.0405
R877 X1.n785 X1.n784 0.0405
R878 X1.n784 X1.n783 0.0405
R879 X1.n783 X1.n776 0.0405
R880 X1.n779 X1.n776 0.0405
R881 X1.n779 X1.n778 0.0405
R882 X1.n778 X1.n428 0.0405
R883 X1.n880 X1.n428 0.0405
R884 X1.n881 X1.n880 0.0405
R885 X1.n883 X1.n881 0.0405
R886 X1.n883 X1.n882 0.0405
R887 X1.n882 X1.n403 0.0405
R888 X1.n933 X1.n403 0.0405
R889 X1.n934 X1.n933 0.0405
R890 X1.n935 X1.n384 0.0405
R891 X1.n976 X1.n384 0.0405
R892 X1.n977 X1.n976 0.0405
R893 X1.n983 X1.n977 0.0405
R894 X1.n983 X1.n982 0.0405
R895 X1.n982 X1.n981 0.0405
R896 X1.n981 X1.n978 0.0405
R897 X1.n978 X1.n350 0.0405
R898 X1.n1068 X1.n350 0.0405
R899 X1.n1069 X1.n1068 0.0405
R900 X1.n1070 X1.n1069 0.0405
R901 X1.n1070 X1.n336 0.0405
R902 X1.n1317 X1.n56 0.0360676
R903 X1.n1319 X1.n1318 0.0360676
R904 X1.n936 X1.n402 0.0360676
R905 X1.n935 X1.n934 0.0360676
R906 X1.n1108 X1.n1107 0.0360676
R907 X1.n1108 X1.n326 0.0360676
R908 X1.n1128 X1.n326 0.0360676
R909 X1.n1129 X1.n1128 0.0360676
R910 X1.n1130 X1.n1129 0.0360676
R911 X1.n1130 X1.n312 0.0360676
R912 X1.n1151 X1.n312 0.0360676
R913 X1.n1152 X1.n1151 0.0360676
R914 X1.n1153 X1.n1152 0.0360676
R915 X1.n1154 X1.n1153 0.0360676
R916 X1.n1154 X1.n300 0.0360676
R917 X1.n1182 X1.n300 0.0360676
R918 X1.n1183 X1.n1182 0.0360676
R919 X1.n1184 X1.n1183 0.0360676
R920 X1.n1185 X1.n1184 0.0360676
R921 X1.n1185 X1.n283 0.0360676
R922 X1.n1206 X1.n283 0.0360676
R923 X1.n1207 X1.n1206 0.0360676
R924 X1.n1208 X1.n1207 0.0360676
R925 X1.n1208 X1.n273 0.0360676
R926 X1.n1229 X1.n273 0.0360676
R927 X1.n1230 X1.n1229 0.0360676
R928 X1.n1231 X1.n1230 0.0360676
R929 X1.n1232 X1.n1231 0.0360676
R930 X1.n1232 X1.n262 0.0360676
R931 X1.n1260 X1.n262 0.0360676
R932 X1.n1261 X1.n1260 0.0360676
R933 X1.n1262 X1.n1261 0.0360676
R934 X1.n1262 X1.n253 0.0360676
R935 X1.n1284 X1.n253 0.0360676
R936 X1.n1285 X1.n1284 0.0360676
R937 X1.n1287 X1.n1285 0.0360676
R938 X1.n1287 X1.n1286 0.0360676
R939 X1.n1109 X1.n335 0.0360676
R940 X1.n1109 X1.n327 0.0360676
R941 X1.n1127 X1.n327 0.0360676
R942 X1.n1127 X1.n325 0.0360676
R943 X1.n1131 X1.n325 0.0360676
R944 X1.n1131 X1.n313 0.0360676
R945 X1.n1150 X1.n313 0.0360676
R946 X1.n1150 X1.n311 0.0360676
R947 X1.n1156 X1.n311 0.0360676
R948 X1.n1156 X1.n1155 0.0360676
R949 X1.n1155 X1.n301 0.0360676
R950 X1.n1181 X1.n301 0.0360676
R951 X1.n1181 X1.n299 0.0360676
R952 X1.n1187 X1.n299 0.0360676
R953 X1.n1187 X1.n1186 0.0360676
R954 X1.n1186 X1.n284 0.0360676
R955 X1.n1205 X1.n284 0.0360676
R956 X1.n1205 X1.n282 0.0360676
R957 X1.n1209 X1.n282 0.0360676
R958 X1.n1209 X1.n274 0.0360676
R959 X1.n1228 X1.n274 0.0360676
R960 X1.n1228 X1.n272 0.0360676
R961 X1.n1234 X1.n272 0.0360676
R962 X1.n1234 X1.n1233 0.0360676
R963 X1.n1233 X1.n263 0.0360676
R964 X1.n1259 X1.n263 0.0360676
R965 X1.n1259 X1.n261 0.0360676
R966 X1.n1263 X1.n261 0.0360676
R967 X1.n1263 X1.n254 0.0360676
R968 X1.n1283 X1.n254 0.0360676
R969 X1.n1283 X1.n252 0.0360676
R970 X1.n1288 X1.n252 0.0360676
R971 X1.n1288 X1.n74 0.0360676
R972 X1.n772 X1.n771 0.0360676
R973 X1.n771 X1.n477 0.0360676
R974 X1.n767 X1.n477 0.0360676
R975 X1.n767 X1.n766 0.0360676
R976 X1.n766 X1.n765 0.0360676
R977 X1.n765 X1.n482 0.0360676
R978 X1.n761 X1.n482 0.0360676
R979 X1.n761 X1.n760 0.0360676
R980 X1.n760 X1.n759 0.0360676
R981 X1.n759 X1.n487 0.0360676
R982 X1.n755 X1.n487 0.0360676
R983 X1.n755 X1.n754 0.0360676
R984 X1.n754 X1.n753 0.0360676
R985 X1.n753 X1.n492 0.0360676
R986 X1.n749 X1.n492 0.0360676
R987 X1.n749 X1.n6 0.0360676
R988 X1.n1374 X1.n6 0.0360676
R989 X1.n1374 X1.n1373 0.0360676
R990 X1.n1373 X1.n1372 0.0360676
R991 X1.n1372 X1.n10 0.0360676
R992 X1.n1368 X1.n10 0.0360676
R993 X1.n1368 X1.n1367 0.0360676
R994 X1.n1367 X1.n1366 0.0360676
R995 X1.n1366 X1.n15 0.0360676
R996 X1.n1362 X1.n15 0.0360676
R997 X1.n1362 X1.n1361 0.0360676
R998 X1.n1361 X1.n1360 0.0360676
R999 X1.n1360 X1.n20 0.0360676
R1000 X1.n1356 X1.n20 0.0360676
R1001 X1.n1356 X1.n1355 0.0360676
R1002 X1.n1355 X1.n1354 0.0360676
R1003 X1.n1354 X1.n25 0.0360676
R1004 X1.n1350 X1.n25 0.0360676
R1005 X1.n770 X1.n473 0.0360676
R1006 X1.n770 X1.n769 0.0360676
R1007 X1.n769 X1.n768 0.0360676
R1008 X1.n768 X1.n478 0.0360676
R1009 X1.n764 X1.n478 0.0360676
R1010 X1.n764 X1.n763 0.0360676
R1011 X1.n763 X1.n762 0.0360676
R1012 X1.n762 X1.n483 0.0360676
R1013 X1.n758 X1.n483 0.0360676
R1014 X1.n758 X1.n757 0.0360676
R1015 X1.n757 X1.n756 0.0360676
R1016 X1.n756 X1.n488 0.0360676
R1017 X1.n752 X1.n488 0.0360676
R1018 X1.n752 X1.n751 0.0360676
R1019 X1.n751 X1.n750 0.0360676
R1020 X1.n750 X1.n4 0.0360676
R1021 X1.n1375 X1.n5 0.0360676
R1022 X1.n1371 X1.n5 0.0360676
R1023 X1.n1371 X1.n1370 0.0360676
R1024 X1.n1370 X1.n1369 0.0360676
R1025 X1.n1369 X1.n11 0.0360676
R1026 X1.n1365 X1.n11 0.0360676
R1027 X1.n1365 X1.n1364 0.0360676
R1028 X1.n1364 X1.n1363 0.0360676
R1029 X1.n1363 X1.n16 0.0360676
R1030 X1.n1359 X1.n16 0.0360676
R1031 X1.n1359 X1.n1358 0.0360676
R1032 X1.n1358 X1.n1357 0.0360676
R1033 X1.n1357 X1.n21 0.0360676
R1034 X1.n1353 X1.n21 0.0360676
R1035 X1.n1353 X1.n1352 0.0360676
R1036 X1.n1352 X1.n1351 0.0360676
R1037 X1.n1349 X1.n28 0.0234189
R1038 X1.n41 X1.n26 0.0234189
R1039 X1.n773 X1.n471 0.0234189
R1040 X1.n775 X1.n774 0.0234189
R1041 X1.n1299 X1.n1298 0.0233108
R1042 X1.n1300 X1.n72 0.0233108
R1043 X1.n1105 X1.n337 0.0233108
R1044 X1.n1106 X1.n336 0.0233108
R1045 X1.n1107 X1.n1106 0.0227703
R1046 X1.n1105 X1.n335 0.0227703
R1047 X1.n773 X1.n772 0.0227703
R1048 X1.n774 X1.n473 0.0227703
R1049 X1.n1376 X1.n1375 0.0219054
R1050 X1.n116 X1.n115 0.0188784
R1051 X1.n120 X1.n119 0.0188784
R1052 X1.n124 X1.n123 0.0188784
R1053 X1.n128 X1.n127 0.0188784
R1054 X1.n133 X1.n132 0.0188784
R1055 X1.n145 X1.n144 0.0188784
R1056 X1.n150 X1.n149 0.0188784
R1057 X1.n157 X1.n101 0.0188784
R1058 X1.n160 X1.n159 0.0188784
R1059 X1.n164 X1.n163 0.0188784
R1060 X1.n169 X1.n167 0.0188784
R1061 X1.n178 X1.n177 0.0188784
R1062 X1.n182 X1.n181 0.0188784
R1063 X1.n186 X1.n185 0.0188784
R1064 X1.n190 X1.n189 0.0188784
R1065 X1.n195 X1.n194 0.0188784
R1066 X1.n198 X1.n197 0.0188784
R1067 X1.n206 X1.n205 0.0188784
R1068 X1.n221 X1.n87 0.0188784
R1069 X1.n224 X1.n223 0.0188784
R1070 X1.n228 X1.n227 0.0188784
R1071 X1.n232 X1.n231 0.0188784
R1072 X1.n234 X1.n83 0.0188784
R1073 X1.n805 X1.n804 0.0188784
R1074 X1.n813 X1.n812 0.0188784
R1075 X1.n822 X1.n821 0.0188784
R1076 X1.n832 X1.n831 0.0188784
R1077 X1.n841 X1.n840 0.0188784
R1078 X1.n856 X1.n430 0.0188784
R1079 X1.n877 X1.n432 0.0188784
R1080 X1.n886 X1.n423 0.0188784
R1081 X1.n425 X1.n420 0.0188784
R1082 X1.n906 X1.n413 0.0188784
R1083 X1.n909 X1.n908 0.0188784
R1084 X1.n930 X1.n406 0.0188784
R1085 X1.n939 X1.n938 0.0188784
R1086 X1.n952 X1.n395 0.0188784
R1087 X1.n954 X1.n386 0.0188784
R1088 X1.n973 X1.n388 0.0188784
R1089 X1.n986 X1.n381 0.0188784
R1090 X1.n1000 X1.n375 0.0188784
R1091 X1.n1017 X1.n1016 0.0188784
R1092 X1.n1027 X1.n1025 0.0188784
R1093 X1.n358 X1.n352 0.0188784
R1094 X1.n1065 X1.n353 0.0188784
R1095 X1.n1043 X1.n1042 0.0188784
R1096 X1.n1104 X1.n339 0.0188784
R1097 X1.n1094 X1.n334 0.0188784
R1098 X1.n1114 X1.n1111 0.0188784
R1099 X1.n1112 X1.n328 0.0188784
R1100 X1.n1197 X1.n285 0.0188784
R1101 X1.n1203 X1.n286 0.0188784
R1102 X1.n291 X1.n281 0.0188784
R1103 X1.n1213 X1.n1211 0.0188784
R1104 X1.n548 X1.n474 0.0188784
R1105 X1.n552 X1.n551 0.0188784
R1106 X1.n565 X1.n560 0.0188784
R1107 X1.n563 X1.n562 0.0188784
R1108 X1.n740 X1.n739 0.0188784
R1109 X1.n735 X1.n734 0.0188784
R1110 X1.n730 X1.n729 0.0188784
R1111 X1.n726 X1.n725 0.0188784
R1112 X1.n1341 X1.n38 0.0187703
R1113 X1.n115 X1.n39 0.0187703
R1114 X1.n136 X1.n135 0.0187703
R1115 X1.n144 X1.n143 0.0187703
R1116 X1.n169 X1.n168 0.0187703
R1117 X1.n207 X1.n206 0.0187703
R1118 X1.n212 X1.n211 0.0187703
R1119 X1.n239 X1.n83 0.0187703
R1120 X1.n242 X1.n241 0.0187703
R1121 X1.n789 X1.n788 0.0187703
R1122 X1.n804 X1.n463 0.0187703
R1123 X1.n848 X1.n847 0.0187703
R1124 X1.n856 X1.n855 0.0187703
R1125 X1.n908 X1.n405 0.0187703
R1126 X1.n1001 X1.n1000 0.0187703
R1127 X1.n1009 X1.n1008 0.0187703
R1128 X1.n1043 X1.n348 0.0187703
R1129 X1.n1075 X1.n1074 0.0187703
R1130 X1.n1122 X1.n324 0.0187703
R1131 X1.n1136 X1.n1133 0.0187703
R1132 X1.n1134 X1.n314 0.0187703
R1133 X1.n1148 X1.n315 0.0187703
R1134 X1.n318 X1.n310 0.0187703
R1135 X1.n1159 X1.n1158 0.0187703
R1136 X1.n1164 X1.n1163 0.0187703
R1137 X1.n1166 X1.n302 0.0187703
R1138 X1.n1179 X1.n303 0.0187703
R1139 X1.n1171 X1.n298 0.0187703
R1140 X1.n1190 X1.n1189 0.0187703
R1141 X1.n1195 X1.n1194 0.0187703
R1142 X1.n1226 X1.n276 0.0187703
R1143 X1.n1218 X1.n271 0.0187703
R1144 X1.n1237 X1.n1236 0.0187703
R1145 X1.n1242 X1.n1241 0.0187703
R1146 X1.n1244 X1.n264 0.0187703
R1147 X1.n1257 X1.n265 0.0187703
R1148 X1.n1253 X1.n260 0.0187703
R1149 X1.n1268 X1.n1265 0.0187703
R1150 X1.n1266 X1.n255 0.0187703
R1151 X1.n1281 X1.n256 0.0187703
R1152 X1.n1276 X1.n251 0.0187703
R1153 X1.n1291 X1.n1290 0.0187703
R1154 X1.n576 X1.n575 0.0187703
R1155 X1.n572 X1.n571 0.0187703
R1156 X1.n585 X1.n584 0.0187703
R1157 X1.n590 X1.n589 0.0187703
R1158 X1.n594 X1.n593 0.0187703
R1159 X1.n511 X1.n510 0.0187703
R1160 X1.n604 X1.n603 0.0187703
R1161 X1.n608 X1.n607 0.0187703
R1162 X1.n612 X1.n611 0.0187703
R1163 X1.n617 X1.n616 0.0187703
R1164 X1.n619 X1.n493 0.0187703
R1165 X1.n747 X1.n494 0.0187703
R1166 X1.n715 X1.n714 0.0187703
R1167 X1.n711 X1.n710 0.0187703
R1168 X1.n706 X1.n705 0.0187703
R1169 X1.n701 X1.n700 0.0187703
R1170 X1.n642 X1.n641 0.0187703
R1171 X1.n648 X1.n647 0.0187703
R1172 X1.n688 X1.n686 0.0187703
R1173 X1.n691 X1.n690 0.0187703
R1174 X1.n683 X1.n682 0.0187703
R1175 X1.n661 X1.n660 0.0187703
R1176 X1.n673 X1.n672 0.0187703
R1177 X1.n670 X1.n665 0.0187703
R1178 X1.n119 X1.n112 0.0185541
R1179 X1.n232 X1.n70 0.0185541
R1180 X1.n812 X1.n459 0.0185541
R1181 X1.n1041 X1.n353 0.0185541
R1182 X1.n1125 X1.n329 0.0184459
R1183 X1.n1227 X1.n275 0.0184459
R1184 X1.n522 X1.n480 0.0184459
R1185 X1.n721 X1.n12 0.0184459
R1186 X1.n177 X1.n55 0.0182297
R1187 X1.n931 X1.n930 0.0182297
R1188 X1.n1126 X1.n1125 0.0181216
R1189 X1.n1212 X1.n275 0.0181216
R1190 X1.n522 X1.n479 0.0181216
R1191 X1.n721 X1.n630 0.0181216
R1192 X1.n135 X1.n48 0.0175811
R1193 X1.n211 X1.n64 0.0175811
R1194 X1.n848 X1.n439 0.0175811
R1195 X1.n1008 X1.n371 0.0175811
R1196 X1.n1132 X1.n324 0.0173649
R1197 X1.n1217 X1.n276 0.0173649
R1198 X1.n576 X1.n481 0.0173649
R1199 X1.n715 X1.n13 0.0173649
R1200 X1.n1113 X1.n1112 0.0170405
R1201 X1.n1211 X1.n1210 0.0170405
R1202 X1.n564 X1.n563 0.0170405
R1203 X1.n726 X1.n9 0.0170405
R1204 X1.n149 X1.n49 0.0167162
R1205 X1.n197 X1.n63 0.0167162
R1206 X1.n878 X1.n877 0.0167162
R1207 X1.n986 X1.n985 0.0167162
R1208 X1.n1136 X1.n1135 0.0162838
R1209 X1.n1235 X1.n271 0.0162838
R1210 X1.n571 X1.n516 0.0162838
R1211 X1.n710 X1.n14 0.0162838
R1212 X1.n164 X1.n54 0.0159595
R1213 X1.n185 X1.n58 0.0159595
R1214 X1.n907 X1.n906 0.0159595
R1215 X1.n937 X1.n395 0.0159595
R1216 X1.n1111 X1.n1110 0.0159595
R1217 X1.n291 X1.n290 0.0159595
R1218 X1.n560 X1.n476 0.0159595
R1219 X1.n730 X1.n8 0.0159595
R1220 X1.n1341 X1.n1340 0.0157432
R1221 X1.n241 X1.n240 0.0157432
R1222 X1.n788 X1.n787 0.0157432
R1223 X1.n1075 X1.n1072 0.0157432
R1224 X1.n123 X1.n43 0.0152027
R1225 X1.n228 X1.n69 0.0152027
R1226 X1.n821 X1.n455 0.0152027
R1227 X1.n1066 X1.n352 0.0152027
R1228 X1.n1149 X1.n314 0.0152027
R1229 X1.n1237 X1.n269 0.0152027
R1230 X1.n585 X1.n484 0.0152027
R1231 X1.n705 X1.n638 0.0152027
R1232 X1.n181 X1.n96 0.0148784
R1233 X1.n939 X1.n401 0.0148784
R1234 X1.n1094 X1.n1093 0.0148784
R1235 X1.n1204 X1.n1203 0.0148784
R1236 X1.n552 X1.n475 0.0148784
R1237 X1.n735 X1.n7 0.0148784
R1238 X1.n1376 X1.n4 0.0146622
R1239 X1.n134 X1.n133 0.0141216
R1240 X1.n87 X1.n65 0.0141216
R1241 X1.n841 X1.n443 0.0141216
R1242 X1.n1016 X1.n366 0.0141216
R1243 X1.n317 X1.n315 0.0141216
R1244 X1.n1243 X1.n1242 0.0141216
R1245 X1.n590 X1.n485 0.0141216
R1246 X1.n700 X1.n17 0.0141216
R1247 X1.n1286 X1.n72 0.0137973
R1248 X1.n1298 X1.n74 0.0137973
R1249 X1.n1197 X1.n1196 0.0137973
R1250 X1.n1297 X1.n76 0.0137973
R1251 X1.n739 X1.n738 0.0137973
R1252 X1.n1348 X1.n27 0.0137973
R1253 X1.n1350 X1.n1349 0.0137973
R1254 X1.n1351 X1.n26 0.0137973
R1255 X1.n1295 X1.n1294 0.0134381
R1256 X1.n101 X1.n50 0.0133649
R1257 X1.n196 X1.n195 0.0133649
R1258 X1.n431 X1.n423 0.0133649
R1259 X1.n388 X1.n387 0.0133649
R1260 X1.n1157 X1.n310 0.0130405
R1261 X1.n1258 X1.n264 0.0130405
R1262 X1.n593 X1.n486 0.0130405
R1263 X1.n642 X1.n18 0.0130405
R1264 X1.n1194 X1.n296 0.0128243
R1265 X1.n1291 X1.n1289 0.0128243
R1266 X1.n748 X1.n747 0.0128243
R1267 X1.n671 X1.n670 0.0128243
R1268 X1.n160 X1.n53 0.0126081
R1269 X1.n189 X1.n59 0.0126081
R1270 X1.n426 X1.n425 0.0126081
R1271 X1.n954 X1.n953 0.0126081
R1272 X1.n37 X1.n29 0.0123919
R1273 X1.n75 X1.n73 0.0123919
R1274 X1.n536 X1.n470 0.0123919
R1275 X1.n1073 X1.n338 0.0123919
R1276 X1.n1159 X1.n308 0.0119595
R1277 X1.n1252 X1.n265 0.0119595
R1278 X1.n510 X1.n507 0.0119595
R1279 X1.n648 X1.n19 0.0119595
R1280 X1.n127 X1.n44 0.0118514
R1281 X1.n224 X1.n68 0.0118514
R1282 X1.n831 X1.n451 0.0118514
R1283 X1.n1027 X1.n1026 0.0118514
R1284 X1.n1189 X1.n1188 0.0117432
R1285 X1.n1276 X1.n1275 0.0117432
R1286 X1.n619 X1.n618 0.0117432
R1287 X1.n673 X1.n24 0.0117432
R1288 X1.n1346 X1.n1345 0.0116588
R1289 X1.n1348 X1.n29 0.011527
R1290 X1.n536 X1.n474 0.011527
R1291 X1.n1297 X1.n75 0.0114189
R1292 X1.n1104 X1.n338 0.0114189
R1293 X1.n569 X1.n568 0.0109762
R1294 X1.n581 X1.n580 0.0109762
R1295 X1.n597 X1.n514 0.0109762
R1296 X1.n600 X1.n598 0.0109762
R1297 X1.n599 X1.n500 0.0109762
R1298 X1.n624 X1.n623 0.0109762
R1299 X1.n743 X1.n497 0.0109762
R1300 X1.n632 X1.n631 0.0109762
R1301 X1.n719 X1.n635 0.0109762
R1302 X1.n697 X1.n639 0.0109762
R1303 X1.n696 X1.n695 0.0109762
R1304 X1.n1344 X1.n33 0.0109762
R1305 X1.n110 X1.n33 0.0109762
R1306 X1.n110 X1.n109 0.0109762
R1307 X1.n109 X1.n106 0.0109762
R1308 X1.n139 X1.n106 0.0109762
R1309 X1.n140 X1.n139 0.0109762
R1310 X1.n140 X1.n103 0.0109762
R1311 X1.n153 X1.n103 0.0109762
R1312 X1.n154 X1.n153 0.0109762
R1313 X1.n154 X1.n98 0.0109762
R1314 X1.n172 X1.n98 0.0109762
R1315 X1.n175 X1.n174 0.0109762
R1316 X1.n174 X1.n173 0.0109762
R1317 X1.n173 X1.n92 0.0109762
R1318 X1.n201 X1.n92 0.0109762
R1319 X1.n202 X1.n201 0.0109762
R1320 X1.n202 X1.n89 0.0109762
R1321 X1.n215 X1.n89 0.0109762
R1322 X1.n218 X1.n215 0.0109762
R1323 X1.n218 X1.n217 0.0109762
R1324 X1.n217 X1.n216 0.0109762
R1325 X1.n216 X1.n81 0.0109762
R1326 X1.n245 X1.n81 0.0109762
R1327 X1.n1118 X1.n1117 0.0109762
R1328 X1.n1139 X1.n320 0.0109762
R1329 X1.n1144 X1.n1140 0.0109762
R1330 X1.n1143 X1.n306 0.0109762
R1331 X1.n1176 X1.n1169 0.0109762
R1332 X1.n1175 X1.n294 0.0109762
R1333 X1.n1200 X1.n1199 0.0109762
R1334 X1.n1216 X1.n279 0.0109762
R1335 X1.n1223 X1.n1222 0.0109762
R1336 X1.n1247 X1.n267 0.0109762
R1337 X1.n1248 X1.n258 0.0109762
R1338 X1.n1272 X1.n1271 0.0109762
R1339 X1.n1294 X1.n249 0.0109762
R1340 X1.n568 X1.n525 0.01095
R1341 X1.n580 X1.n569 0.01095
R1342 X1.n581 X1.n514 0.01095
R1343 X1.n598 X1.n597 0.01095
R1344 X1.n600 X1.n599 0.01095
R1345 X1.n623 X1.n500 0.01095
R1346 X1.n743 X1.n624 0.01095
R1347 X1.n631 X1.n497 0.01095
R1348 X1.n719 X1.n632 0.01095
R1349 X1.n639 X1.n635 0.01095
R1350 X1.n697 X1.n696 0.01095
R1351 X1.n695 X1.n694 0.01095
R1352 X1.n175 X1.n172 0.01095
R1353 X1.n246 X1.n245 0.01095
R1354 X1.n1118 X1.n320 0.01095
R1355 X1.n1140 X1.n1139 0.01095
R1356 X1.n1144 X1.n1143 0.01095
R1357 X1.n1169 X1.n306 0.01095
R1358 X1.n1176 X1.n1175 0.01095
R1359 X1.n1199 X1.n294 0.01095
R1360 X1.n1200 X1.n279 0.01095
R1361 X1.n1223 X1.n1216 0.01095
R1362 X1.n1222 X1.n267 0.01095
R1363 X1.n1248 X1.n1247 0.01095
R1364 X1.n1271 X1.n258 0.01095
R1365 X1.n1272 X1.n249 0.01095
R1366 X1.n1165 X1.n1164 0.0108784
R1367 X1.n1264 X1.n260 0.0108784
R1368 X1.n604 X1.n489 0.0108784
R1369 X1.n689 X1.n688 0.0108784
R1370 X1.n128 X1.n45 0.0107703
R1371 X1.n223 X1.n222 0.0107703
R1372 X1.n832 X1.n447 0.0107703
R1373 X1.n1025 X1.n361 0.0107703
R1374 X1.n1171 X1.n1170 0.0106622
R1375 X1.n1282 X1.n1281 0.0106622
R1376 X1.n616 X1.n491 0.0106622
R1377 X1.n660 X1.n23 0.0106622
R1378 X1.n1345 X1.n1344 0.0106095
R1379 X1.n159 X1.n158 0.0100135
R1380 X1.n190 X1.n60 0.0100135
R1381 X1.n885 X1.n420 0.0100135
R1382 X1.n974 X1.n386 0.0100135
R1383 X1.n1180 X1.n302 0.0097973
R1384 X1.n1268 X1.n1267 0.0097973
R1385 X1.n608 X1.n490 0.0097973
R1386 X1.n691 X1.n22 0.0097973
R1387 X1.n1346 X1.n32 0.00967266
R1388 X1.n1180 X1.n1179 0.00958108
R1389 X1.n1267 X1.n1266 0.00958108
R1390 X1.n611 X1.n490 0.00958108
R1391 X1.n683 X1.n22 0.00958108
R1392 X1.n158 X1.n157 0.00925676
R1393 X1.n194 X1.n60 0.00925676
R1394 X1.n886 X1.n885 0.00925676
R1395 X1.n974 X1.n973 0.00925676
R1396 X1.n623 X1.n499 0.00880612
R1397 X1.n1170 X1.n303 0.00871622
R1398 X1.n1282 X1.n255 0.00871622
R1399 X1.n612 X1.n491 0.00871622
R1400 X1.n682 X1.n23 0.00871622
R1401 X1.n132 X1.n45 0.0085
R1402 X1.n222 X1.n221 0.0085
R1403 X1.n840 X1.n447 0.0085
R1404 X1.n1017 X1.n361 0.0085
R1405 X1.n1166 X1.n1165 0.0085
R1406 X1.n1265 X1.n1264 0.0085
R1407 X1.n607 X1.n489 0.0085
R1408 X1.n690 X1.n689 0.0085
R1409 X1.n1117 X1.n331 0.00809524
R1410 X1.n666 X1.n663 0.00778095
R1411 X1.n1188 X1.n298 0.00763514
R1412 X1.n1275 X1.n256 0.00763514
R1413 X1.n618 X1.n617 0.00763514
R1414 X1.n661 X1.n24 0.00763514
R1415 X1.n124 X1.n44 0.00741892
R1416 X1.n227 X1.n68 0.00741892
R1417 X1.n822 X1.n451 0.00741892
R1418 X1.n1026 X1.n358 0.00741892
R1419 X1.n1163 X1.n308 0.00741892
R1420 X1.n1253 X1.n1252 0.00741892
R1421 X1.n603 X1.n507 0.00741892
R1422 X1.n686 X1.n19 0.00741892
R1423 X1.n694 X1.n652 0.00725714
R1424 X1.n666 X1.n32 0.00707381
R1425 X1.n38 X1.n37 0.00698649
R1426 X1.n242 X1.n73 0.00698649
R1427 X1.n789 X1.n470 0.00698649
R1428 X1.n1074 X1.n1073 0.00698649
R1429 X1.n546 X1.n525 0.00696162
R1430 X1.n246 X1.n80 0.00691667
R1431 X1.n163 X1.n53 0.00666216
R1432 X1.n186 X1.n59 0.00666216
R1433 X1.n426 X1.n413 0.00666216
R1434 X1.n953 X1.n952 0.00666216
R1435 X1.n1190 X1.n296 0.00655405
R1436 X1.n1289 X1.n251 0.00655405
R1437 X1.n748 X1.n493 0.00655405
R1438 X1.n672 X1.n671 0.00655405
R1439 X1.n1158 X1.n1157 0.00633784
R1440 X1.n1258 X1.n1257 0.00633784
R1441 X1.n511 X1.n486 0.00633784
R1442 X1.n647 X1.n18 0.00633784
R1443 X1.n150 X1.n50 0.00590541
R1444 X1.n198 X1.n196 0.00590541
R1445 X1.n432 X1.n431 0.00590541
R1446 X1.n387 X1.n381 0.00590541
R1447 X1.n627 X1.n497 0.00588776
R1448 X1.n556 X1.n525 0.00588776
R1449 X1.n1196 X1.n1195 0.00547297
R1450 X1.n1290 X1.n76 0.00547297
R1451 X1.n738 X1.n494 0.00547297
R1452 X1.n665 X1.n27 0.00547297
R1453 X1.n318 X1.n317 0.00525676
R1454 X1.n1244 X1.n1243 0.00525676
R1455 X1.n594 X1.n485 0.00525676
R1456 X1.n641 X1.n17 0.00525676
R1457 X1.n136 X1.n134 0.00514865
R1458 X1.n212 X1.n65 0.00514865
R1459 X1.n847 X1.n443 0.00514865
R1460 X1.n1009 X1.n366 0.00514865
R1461 X1.n1295 X1.n248 0.00440238
R1462 X1.n178 X1.n96 0.00439189
R1463 X1.n406 X1.n401 0.00439189
R1464 X1.n1093 X1.n339 0.00439189
R1465 X1.n1204 X1.n285 0.00439189
R1466 X1.n548 X1.n475 0.00439189
R1467 X1.n740 X1.n7 0.00439189
R1468 X1.n35 X1.n34 0.00425921
R1469 X1.n1342 X1.n36 0.00425921
R1470 X1.n129 X1.n126 0.00425921
R1471 X1.n131 X1.n107 0.00425921
R1472 X1.n146 X1.n104 0.00425921
R1473 X1.n151 X1.n148 0.00425921
R1474 X1.n156 X1.n102 0.00425921
R1475 X1.n161 X1.n100 0.00425921
R1476 X1.n179 X1.n176 0.00425921
R1477 X1.n191 X1.n188 0.00425921
R1478 X1.n193 X1.n93 0.00425921
R1479 X1.n199 X1.n91 0.00425921
R1480 X1.n204 X1.n90 0.00425921
R1481 X1.n220 X1.n88 0.00425921
R1482 X1.n225 X1.n86 0.00425921
R1483 X1.n238 X1.n82 0.00425921
R1484 X1.n243 X1.n77 0.00425921
R1485 X1.n333 X1.n330 0.00425921
R1486 X1.n1124 X1.n1123 0.00425921
R1487 X1.n1120 X1.n321 0.00425921
R1488 X1.n1137 X1.n323 0.00425921
R1489 X1.n1162 X1.n1160 0.00425921
R1490 X1.n1167 X1.n307 0.00425921
R1491 X1.n1178 X1.n304 0.00425921
R1492 X1.n1172 X1.n305 0.00425921
R1493 X1.n1198 X1.n287 0.00425921
R1494 X1.n1214 X1.n280 0.00425921
R1495 X1.n1225 X1.n277 0.00425921
R1496 X1.n1219 X1.n278 0.00425921
R1497 X1.n1220 X1.n270 0.00425921
R1498 X1.n1255 X1.n1254 0.00425921
R1499 X1.n1250 X1.n259 0.00425921
R1500 X1.n1269 X1.n257 0.00425921
R1501 X1.n1280 X1.n1274 0.00425921
R1502 X1.n606 X1.n605 0.00425921
R1503 X1.n610 X1.n609 0.00425921
R1504 X1.n687 X1.n653 0.00425921
R1505 X1.n692 X1.n684 0.00425921
R1506 X1.n679 X1.n657 0.00424524
R1507 X1.n114 X1.n36 0.0042371
R1508 X1.n118 X1.n117 0.0042371
R1509 X1.n122 X1.n121 0.0042371
R1510 X1.n126 X1.n125 0.0042371
R1511 X1.n137 X1.n105 0.0042371
R1512 X1.n142 X1.n104 0.0042371
R1513 X1.n162 X1.n161 0.0042371
R1514 X1.n166 X1.n165 0.0042371
R1515 X1.n170 X1.n97 0.0042371
R1516 X1.n176 X1.n97 0.0042371
R1517 X1.n180 X1.n179 0.0042371
R1518 X1.n184 X1.n183 0.0042371
R1519 X1.n188 X1.n187 0.0042371
R1520 X1.n208 X1.n90 0.0042371
R1521 X1.n213 X1.n210 0.0042371
R1522 X1.n226 X1.n225 0.0042371
R1523 X1.n230 X1.n229 0.0042371
R1524 X1.n235 X1.n233 0.0042371
R1525 X1.n238 X1.n237 0.0042371
R1526 X1.n1096 X1.n332 0.0042371
R1527 X1.n1115 X1.n333 0.0042371
R1528 X1.n323 X1.n322 0.0042371
R1529 X1.n1147 X1.n1146 0.0042371
R1530 X1.n1141 X1.n319 0.0042371
R1531 X1.n1160 X1.n309 0.0042371
R1532 X1.n1173 X1.n1172 0.0042371
R1533 X1.n1191 X1.n297 0.0042371
R1534 X1.n1193 X1.n295 0.0042371
R1535 X1.n1198 X1.n295 0.0042371
R1536 X1.n1202 X1.n287 0.0042371
R1537 X1.n293 X1.n292 0.0042371
R1538 X1.n288 X1.n280 0.0042371
R1539 X1.n1238 X1.n270 0.0042371
R1540 X1.n1240 X1.n268 0.0042371
R1541 X1.n1245 X1.n266 0.0042371
R1542 X1.n1256 X1.n1255 0.0042371
R1543 X1.n1280 X1.n1279 0.0042371
R1544 X1.n1277 X1.n250 0.0042371
R1545 X1.n1292 X1.n78 0.0042371
R1546 X1.n1296 X1.n78 0.0042371
R1547 X1.n566 X1.n559 0.0042371
R1548 X1.n591 X1.n588 0.0042371
R1549 X1.n595 X1.n592 0.0042371
R1550 X1.n746 X1.n745 0.0042371
R1551 X1.n728 X1.n727 0.0042371
R1552 X1.n702 X1.n699 0.0042371
R1553 X1.n643 X1.n640 0.0042371
R1554 X1.n674 X1.n664 0.0042371
R1555 X1.n669 X1.n668 0.0042371
R1556 X1.n1102 X1.n1101 0.00423273
R1557 X1.n745 X1.n744 0.00423268
R1558 X1.n1090 X1.n1089 0.00422178
R1559 X1.n531 X1.n528 0.00422178
R1560 X1.n656 X1.n652 0.00421905
R1561 X1.n1149 X1.n1148 0.00417568
R1562 X1.n1241 X1.n269 0.00417568
R1563 X1.n589 X1.n484 0.00417568
R1564 X1.n701 X1.n638 0.00417568
R1565 X1.n117 X1.n113 0.00410442
R1566 X1.n236 X1.n235 0.00410442
R1567 X1.n120 X1.n43 0.00406757
R1568 X1.n231 X1.n69 0.00406757
R1569 X1.n813 X1.n455 0.00406757
R1570 X1.n1066 X1.n1065 0.00406757
R1571 X1.n503 X1.n502 0.00402269
R1572 X1.n523 X1.n519 0.00398793
R1573 X1.n722 X1.n720 0.00398793
R1574 X1.n1124 X1.n1119 0.00397174
R1575 X1.n1178 X1.n1177 0.00397174
R1576 X1.n1215 X1.n277 0.00397174
R1577 X1.n1273 X1.n257 0.00397174
R1578 X1.n156 X1.n155 0.00394963
R1579 X1.n193 X1.n192 0.00394963
R1580 X1.n558 X1.n557 0.00394626
R1581 X1.n732 X1.n731 0.00394626
R1582 X1.n550 X1.n549 0.00393696
R1583 X1.n741 X1.n737 0.00393696
R1584 X1.n574 X1.n573 0.00390294
R1585 X1.n713 X1.n712 0.00390294
R1586 X1.n615 X1.n498 0.00389381
R1587 X1.n583 X1.n582 0.00385851
R1588 X1.n601 X1.n508 0.00385851
R1589 X1.n708 X1.n707 0.00385851
R1590 X1.n650 X1.n649 0.00385851
R1591 X1.n583 X1.n515 0.00380768
R1592 X1.n707 X1.n637 0.00380768
R1593 X1.n513 X1.n508 0.00380053
R1594 X1.n649 X1.n645 0.00380053
R1595 X1.n131 X1.n130 0.00379484
R1596 X1.n220 X1.n219 0.00379484
R1597 X1.n1103 X1.n342 0.00379484
R1598 X1.n1347 X1.n31 0.00377273
R1599 X1.n559 X1.n521 0.0037725
R1600 X1.n615 X1.n614 0.0037725
R1601 X1.n727 X1.n629 0.0037725
R1602 X1.n678 X1.n677 0.00374762
R1603 X1.n1147 X1.n316 0.0037285
R1604 X1.n1240 X1.n1239 0.0037285
R1605 X1.n1142 X1.n1141 0.00370639
R1606 X1.n1249 X1.n266 0.00370639
R1607 X1.n676 X1.n663 0.00369524
R1608 X1.n141 X1.n105 0.00366216
R1609 X1.n210 X1.n209 0.00366216
R1610 X1.n681 X1.n680 0.00366216
R1611 X1.n655 X1.n654 0.00364005
R1612 X1.n1340 X1.n39 0.00363514
R1613 X1.n240 X1.n239 0.00363514
R1614 X1.n787 X1.n463 0.00363514
R1615 X1.n1072 X1.n348 0.00363514
R1616 X1.n1100 X1.n1099 0.00359048
R1617 X1.n610 X1.n504 0.00358532
R1618 X1.n742 X1.n496 0.00358218
R1619 X1.n532 X1.n531 0.00357902
R1620 X1.n1089 X1.n343 0.00357902
R1621 X1.n524 X1.n523 0.00357098
R1622 X1.n723 X1.n722 0.00357098
R1623 X1.n148 X1.n147 0.00348526
R1624 X1.n203 X1.n91 0.00348526
R1625 X1.n588 X1.n587 0.003457
R1626 X1.n703 X1.n702 0.003457
R1627 X1.n592 X1.n509 0.00344926
R1628 X1.n644 X1.n643 0.00344926
R1629 X1.n1138 X1.n321 0.00344103
R1630 X1.n1161 X1.n307 0.00344103
R1631 X1.n1221 X1.n1219 0.00344103
R1632 X1.n1251 X1.n1250 0.00344103
R1633 X1.n602 X1.n506 0.00343273
R1634 X1.n685 X1.n651 0.00343273
R1635 X1.n518 X1.n517 0.00341839
R1636 X1.n709 X1.n636 0.00341839
R1637 X1.n719 X1.n634 0.00341837
R1638 X1.n580 X1.n520 0.00341837
R1639 X1.n1098 X1.n331 0.00335476
R1640 X1.n122 X1.n108 0.00335258
R1641 X1.n229 X1.n85 0.00335258
R1642 X1.n573 X1.n518 0.0033136
R1643 X1.n712 X1.n636 0.0033136
R1644 X1.n167 X1.n54 0.00331081
R1645 X1.n182 X1.n58 0.00331081
R1646 X1.n909 X1.n907 0.00331081
R1647 X1.n938 X1.n937 0.00331081
R1648 X1.n1110 X1.n334 0.00331081
R1649 X1.n290 X1.n286 0.00331081
R1650 X1.n551 X1.n476 0.00331081
R1651 X1.n734 X1.n8 0.00331081
R1652 X1.n512 X1.n509 0.00330444
R1653 X1.n646 X1.n644 0.00330444
R1654 X1.n605 X1.n506 0.0032992
R1655 X1.n687 X1.n651 0.0032992
R1656 X1.n587 X1.n586 0.00329663
R1657 X1.n704 X1.n703 0.00329663
R1658 X1.n662 X1.n659 0.00324201
R1659 X1.n165 X1.n99 0.00319779
R1660 X1.n184 X1.n94 0.00319779
R1661 X1.n1174 X1.n297 0.00319779
R1662 X1.n1278 X1.n1277 0.00319779
R1663 X1.n675 X1.n674 0.00319779
R1664 X1.n1116 X1.n332 0.00317568
R1665 X1.n292 X1.n289 0.00317568
R1666 X1.n567 X1.n558 0.00317568
R1667 X1.n731 X1.n628 0.00317568
R1668 X1.n561 X1.n524 0.00316007
R1669 X1.n724 X1.n723 0.00316007
R1670 X1.n613 X1.n504 0.00314581
R1671 X1.n1095 X1.n1092 0.00310934
R1672 X1.n1135 X1.n1134 0.00309459
R1673 X1.n1236 X1.n1235 0.00309459
R1674 X1.n584 X1.n516 0.00309459
R1675 X1.n706 X1.n14 0.00309459
R1676 X1.n1343 X1.n35 0.003043
R1677 X1.n244 X1.n243 0.003043
R1678 X1.n818 X1.n816 0.0029881
R1679 X1.n851 X1.n441 0.0029881
R1680 X1.n874 X1.n866 0.0029881
R1681 X1.n990 X1.n989 0.0029881
R1682 X1.n561 X1.n521 0.00298054
R1683 X1.n614 X1.n613 0.00298054
R1684 X1.n724 X1.n629 0.00298054
R1685 X1.n1005 X1.n369 0.0029619
R1686 X1.n1037 X1.n1036 0.0029619
R1687 X1.n513 X1.n512 0.00293083
R1688 X1.n646 X1.n645 0.00293083
R1689 X1.n586 X1.n515 0.0029237
R1690 X1.n704 X1.n637 0.0029237
R1691 X1.n171 X1.n166 0.00291032
R1692 X1.n183 X1.n95 0.00291032
R1693 X1.n1097 X1.n1096 0.00291032
R1694 X1.n1192 X1.n1191 0.00291032
R1695 X1.n1201 X1.n293 0.00291032
R1696 X1.n1293 X1.n250 0.00291032
R1697 X1.n502 X1.n495 0.00291032
R1698 X1.n667 X1.n664 0.00291032
R1699 X1.n582 X1.n517 0.00289527
R1700 X1.n602 X1.n601 0.00289527
R1701 X1.n709 X1.n708 0.00289527
R1702 X1.n685 X1.n650 0.00289527
R1703 X1.n533 X1.n532 0.00287188
R1704 X1.n1087 X1.n343 0.00284569
R1705 X1.n501 X1.n498 0.00283826
R1706 X1.n248 X1.n80 0.00283095
R1707 X1.n553 X1.n550 0.00279542
R1708 X1.n737 X1.n736 0.00279542
R1709 X1.n570 X1.n519 0.00276679
R1710 X1.n720 X1.n633 0.00276679
R1711 X1.n121 X1.n111 0.00275553
R1712 X1.n230 X1.n84 0.00275553
R1713 X1.n34 X1.n30 0.00273342
R1714 X1.n1296 X1.n77 0.00273342
R1715 X1.n541 X1.n533 0.00272619
R1716 X1.n541 X1.n540 0.00272619
R1717 X1.n792 X1.n468 0.00272619
R1718 X1.n794 X1.n793 0.00272619
R1719 X1.n802 X1.n801 0.00272619
R1720 X1.n810 X1.n457 0.00272619
R1721 X1.n815 X1.n457 0.00272619
R1722 X1.n817 X1.n453 0.00272619
R1723 X1.n825 X1.n453 0.00272619
R1724 X1.n827 X1.n449 0.00272619
R1725 X1.n835 X1.n449 0.00272619
R1726 X1.n843 X1.n445 0.00272619
R1727 X1.n844 X1.n843 0.00272619
R1728 X1.n853 X1.n852 0.00272619
R1729 X1.n853 X1.n437 0.00272619
R1730 X1.n861 X1.n435 0.00272619
R1731 X1.n865 X1.n435 0.00272619
R1732 X1.n873 X1.n872 0.00272619
R1733 X1.n868 X1.n867 0.00272619
R1734 X1.n891 X1.n418 0.00272619
R1735 X1.n901 X1.n900 0.00272619
R1736 X1.n904 X1.n901 0.00272619
R1737 X1.n912 X1.n411 0.00272619
R1738 X1.n913 X1.n912 0.00272619
R1739 X1.n914 X1.n913 0.00272619
R1740 X1.n928 X1.n927 0.00272619
R1741 X1.n942 X1.n399 0.00272619
R1742 X1.n943 X1.n942 0.00272619
R1743 X1.n949 X1.n948 0.00272619
R1744 X1.n950 X1.n949 0.00272619
R1745 X1.n950 X1.n393 0.00272619
R1746 X1.n959 X1.n391 0.00272619
R1747 X1.n963 X1.n391 0.00272619
R1748 X1.n969 X1.n968 0.00272619
R1749 X1.n968 X1.n965 0.00272619
R1750 X1.n995 X1.n377 0.00272619
R1751 X1.n1004 X1.n1003 0.00272619
R1752 X1.n1012 X1.n1011 0.00272619
R1753 X1.n1014 X1.n1013 0.00272619
R1754 X1.n1023 X1.n1022 0.00272619
R1755 X1.n1032 X1.n356 0.00272619
R1756 X1.n1036 X1.n356 0.00272619
R1757 X1.n1063 X1.n1062 0.00272619
R1758 X1.n1062 X1.n1061 0.00272619
R1759 X1.n1061 X1.n1038 0.00272619
R1760 X1.n1052 X1.n1040 0.00272619
R1761 X1.n1052 X1.n1051 0.00272619
R1762 X1.n1045 X1.n346 0.00272619
R1763 X1.n1078 X1.n346 0.00272619
R1764 X1.n1085 X1.n1084 0.00272619
R1765 X1.n1087 X1.n1086 0.00272619
R1766 X1.n540 X1.n539 0.0027
R1767 X1.n793 X1.n792 0.0027
R1768 X1.n802 X1.n800 0.0027
R1769 X1.n810 X1.n809 0.0027
R1770 X1.n818 X1.n817 0.0027
R1771 X1.n845 X1.n844 0.0027
R1772 X1.n872 X1.n867 0.0027
R1773 X1.n891 X1.n890 0.0027
R1774 X1.n900 X1.n416 0.0027
R1775 X1.n928 X1.n920 0.0027
R1776 X1.n921 X1.n399 0.0027
R1777 X1.n965 X1.n379 0.0027
R1778 X1.n991 X1.n377 0.0027
R1779 X1.n1003 X1.n373 0.0027
R1780 X1.n1014 X1.n1012 0.0027
R1781 X1.n1023 X1.n1021 0.0027
R1782 X1.n1032 X1.n1031 0.0027
R1783 X1.n1079 X1.n1078 0.0027
R1784 X1.n1086 X1.n1085 0.0027
R1785 X1.n845 X1.n441 0.00264762
R1786 X1.n1011 X1.n369 0.00264762
R1787 X1.n1121 X1.n1120 0.00264496
R1788 X1.n1224 X1.n278 0.00264496
R1789 X1.n1168 X1.n1167 0.00262285
R1790 X1.n1270 X1.n259 0.00262285
R1791 X1.n606 X1.n505 0.00262285
R1792 X1.n693 X1.n653 0.00262285
R1793 X1.n866 X1.n865 0.00262143
R1794 X1.n991 X1.n990 0.00262143
R1795 X1.n152 X1.n151 0.00260074
R1796 X1.n200 X1.n199 0.00260074
R1797 X1.n820 X1.n456 0.00257862
R1798 X1.n1035 X1.n354 0.00257862
R1799 X1.n989 X1.n379 0.00256905
R1800 X1.n145 X1.n49 0.00255405
R1801 X1.n205 X1.n63 0.00255405
R1802 X1.n878 X1.n430 0.00255405
R1803 X1.n985 X1.n375 0.00255405
R1804 X1.n874 X1.n873 0.00254286
R1805 X1.n1005 X1.n1004 0.00254286
R1806 X1.n876 X1.n875 0.0025344
R1807 X1.n852 X1.n851 0.00251667
R1808 X1.n988 X1.n987 0.00251228
R1809 X1.n744 X1.n496 0.00249519
R1810 X1.n545 X1.n544 0.0024936
R1811 X1.n816 X1.n815 0.00246429
R1812 X1.n1063 X1.n1037 0.00246429
R1813 X1.n138 X1.n137 0.00244595
R1814 X1.n214 X1.n213 0.00244595
R1815 X1.n836 X1.n835 0.0024381
R1816 X1.n1021 X1.n1020 0.0024381
R1817 X1.n849 X1.n442 0.00242383
R1818 X1.n1007 X1.n370 0.00242383
R1819 X1.n679 X1.n678 0.00238571
R1820 X1.n1101 X1.n1100 0.00238571
R1821 X1.n799 X1.n466 0.00238571
R1822 X1.n808 X1.n461 0.00238571
R1823 X1.n828 X1.n826 0.00238571
R1824 X1.n837 X1.n836 0.00238571
R1825 X1.n860 X1.n859 0.00238571
R1826 X1.n889 X1.n421 0.00238571
R1827 X1.n896 X1.n895 0.00238571
R1828 X1.n919 X1.n409 0.00238571
R1829 X1.n926 X1.n922 0.00238571
R1830 X1.n944 X1.n943 0.00238571
R1831 X1.n958 X1.n957 0.00238571
R1832 X1.n970 X1.n964 0.00238571
R1833 X1.n997 X1.n996 0.00238571
R1834 X1.n1020 X1.n364 0.00238571
R1835 X1.n1030 X1.n359 0.00238571
R1836 X1.n1057 X1.n1056 0.00238571
R1837 X1.n1050 X1.n1046 0.00238571
R1838 X1.n791 X1.n790 0.00237961
R1839 X1.n795 X1.n467 0.00237961
R1840 X1.n803 X1.n465 0.00237961
R1841 X1.n811 X1.n458 0.00237961
R1842 X1.n814 X1.n458 0.00237961
R1843 X1.n823 X1.n454 0.00237961
R1844 X1.n824 X1.n823 0.00237961
R1845 X1.n833 X1.n450 0.00237961
R1846 X1.n834 X1.n833 0.00237961
R1847 X1.n842 X1.n446 0.00237961
R1848 X1.n842 X1.n444 0.00237961
R1849 X1.n854 X1.n440 0.00237961
R1850 X1.n854 X1.n438 0.00237961
R1851 X1.n863 X1.n862 0.00237961
R1852 X1.n864 X1.n863 0.00237961
R1853 X1.n871 X1.n434 0.00237961
R1854 X1.n870 X1.n869 0.00237961
R1855 X1.n893 X1.n892 0.00237961
R1856 X1.n899 X1.n414 0.00237961
R1857 X1.n905 X1.n414 0.00237961
R1858 X1.n911 X1.n910 0.00237961
R1859 X1.n911 X1.n410 0.00237961
R1860 X1.n915 X1.n410 0.00237961
R1861 X1.n929 X1.n408 0.00237961
R1862 X1.n941 X1.n940 0.00237961
R1863 X1.n941 X1.n398 0.00237961
R1864 X1.n947 X1.n396 0.00237961
R1865 X1.n951 X1.n396 0.00237961
R1866 X1.n951 X1.n394 0.00237961
R1867 X1.n961 X1.n960 0.00237961
R1868 X1.n962 X1.n961 0.00237961
R1869 X1.n967 X1.n390 0.00237961
R1870 X1.n967 X1.n966 0.00237961
R1871 X1.n994 X1.n993 0.00237961
R1872 X1.n1002 X1.n372 0.00237961
R1873 X1.n1010 X1.n367 0.00237961
R1874 X1.n1015 X1.n368 0.00237961
R1875 X1.n1024 X1.n363 0.00237961
R1876 X1.n1034 X1.n1033 0.00237961
R1877 X1.n1035 X1.n1034 0.00237961
R1878 X1.n1064 X1.n355 0.00237961
R1879 X1.n1060 X1.n355 0.00237961
R1880 X1.n1060 X1.n1059 0.00237961
R1881 X1.n1054 X1.n1053 0.00237961
R1882 X1.n1053 X1.n1044 0.00237961
R1883 X1.n1076 X1.n347 0.00237961
R1884 X1.n1077 X1.n1076 0.00237961
R1885 X1.n1083 X1.n340 0.00237961
R1886 X1.n1146 X1.n1145 0.00237961
R1887 X1.n1145 X1.n319 0.00237961
R1888 X1.n1246 X1.n268 0.00237961
R1889 X1.n1246 X1.n1245 0.00237961
R1890 X1.n543 X1.n527 0.00237961
R1891 X1.n555 X1.n526 0.00237961
R1892 X1.n596 X1.n591 0.00237961
R1893 X1.n596 X1.n595 0.00237961
R1894 X1.n621 X1.n620 0.00237961
R1895 X1.n733 X1.n626 0.00237961
R1896 X1.n699 X1.n698 0.00237961
R1897 X1.n698 X1.n640 0.00237961
R1898 X1.n890 X1.n889 0.00235952
R1899 X1.n902 X1.n411 0.00235952
R1900 X1.n538 X1.n529 0.00235749
R1901 X1.n791 X1.n467 0.00235749
R1902 X1.n803 X1.n464 0.00235749
R1903 X1.n811 X1.n460 0.00235749
R1904 X1.n819 X1.n454 0.00235749
R1905 X1.n846 X1.n444 0.00235749
R1906 X1.n871 X1.n870 0.00235749
R1907 X1.n892 X1.n419 0.00235749
R1908 X1.n899 X1.n898 0.00235749
R1909 X1.n929 X1.n407 0.00235749
R1910 X1.n940 X1.n400 0.00235749
R1911 X1.n966 X1.n380 0.00235749
R1912 X1.n993 X1.n992 0.00235749
R1913 X1.n1002 X1.n374 0.00235749
R1914 X1.n1015 X1.n367 0.00235749
R1915 X1.n1024 X1.n362 0.00235749
R1916 X1.n1033 X1.n357 0.00235749
R1917 X1.n1077 X1.n345 0.00235749
R1918 X1.n578 X1.n577 0.00235749
R1919 X1.n717 X1.n716 0.00235749
R1920 X1.n964 X1.n963 0.00233333
R1921 X1.n846 X1.n442 0.00231327
R1922 X1.n1010 X1.n370 0.00231327
R1923 X1.n539 X1.n535 0.00230714
R1924 X1.n1080 X1.n1079 0.00230714
R1925 X1.n1084 X1.n344 0.00230714
R1926 X1.n138 X1.n107 0.00229115
R1927 X1.n214 X1.n88 0.00229115
R1928 X1.n864 X1.n433 0.00229115
R1929 X1.n992 X1.n378 0.00229115
R1930 X1.n534 X1.n468 0.00228095
R1931 X1.n801 X1.n461 0.00228095
R1932 X1.n1056 X1.n1040 0.00225476
R1933 X1.n988 X1.n380 0.00224693
R1934 X1.n1114 X1.n1113 0.00222973
R1935 X1.n1210 X1.n281 0.00222973
R1936 X1.n565 X1.n564 0.00222973
R1937 X1.n729 X1.n9 0.00222973
R1938 X1.n875 X1.n434 0.00222482
R1939 X1.n1006 X1.n372 0.00222482
R1940 X1.n850 X1.n440 0.0022027
R1941 X1.n904 X1.n903 0.00220238
R1942 X1.n948 X1.n397 0.00220238
R1943 X1.n920 X1.n919 0.00217619
R1944 X1.n927 X1.n926 0.00217619
R1945 X1.n742 X1.n741 0.00217613
R1946 X1.n814 X1.n456 0.00215848
R1947 X1.n1064 X1.n354 0.00215848
R1948 X1.n152 X1.n102 0.00213636
R1949 X1.n200 X1.n93 0.00213636
R1950 X1.n834 X1.n448 0.00213636
R1951 X1.n1019 X1.n362 0.00213636
R1952 X1.n1168 X1.n304 0.00211425
R1953 X1.n1270 X1.n1269 0.00211425
R1954 X1.n609 X1.n505 0.00211425
R1955 X1.n693 X1.n692 0.00211425
R1956 X1.n1099 X1.n1098 0.00209762
R1957 X1.n800 X1.n799 0.00209762
R1958 X1.n945 X1.n398 0.00209214
R1959 X1.n1123 X1.n1121 0.00209214
R1960 X1.n1225 X1.n1224 0.00209214
R1961 X1.n579 X1.n570 0.00209214
R1962 X1.n718 X1.n633 0.00209214
R1963 X1.n1051 X1.n1050 0.00207143
R1964 X1.n888 X1.n419 0.00207002
R1965 X1.n910 X1.n412 0.00207002
R1966 X1.n962 X1.n389 0.00204791
R1967 X1.n538 X1.n537 0.0020258
R1968 X1.n1081 X1.n345 0.0020258
R1969 X1.n1083 X1.n1082 0.0020258
R1970 X1.n895 X1.n418 0.00201905
R1971 X1.n1133 X1.n1132 0.00201351
R1972 X1.n1218 X1.n1217 0.00201351
R1973 X1.n572 X1.n481 0.00201351
R1974 X1.n711 X1.n13 0.00201351
R1975 X1.n118 X1.n111 0.00200369
R1976 X1.n233 X1.n84 0.00200369
R1977 X1.n790 X1.n469 0.00200369
R1978 X1.n465 X1.n462 0.00200369
R1979 X1.n1102 X1.n1090 0.00200107
R1980 X1.n544 X1.n528 0.00200107
R1981 X1.n546 X1.n545 0.00200107
R1982 X1.n959 X1.n958 0.00199286
R1983 X1.n1055 X1.n1054 0.00198157
R1984 X1.n905 X1.n415 0.00193735
R1985 X1.n947 X1.n946 0.00193735
R1986 X1.n918 X1.n407 0.00191523
R1987 X1.n925 X1.n408 0.00191523
R1988 X1.n1103 X1.n341 0.00191523
R1989 X1.n1296 X1.n79 0.00191523
R1990 X1.n543 X1.n542 0.00191523
R1991 X1.n547 X1.n527 0.00191523
R1992 X1.n828 X1.n827 0.00191429
R1993 X1.n1022 X1.n359 0.00191429
R1994 X1.n839 X1.n838 0.00187101
R1995 X1.n577 X1.n574 0.00185493
R1996 X1.n716 X1.n713 0.00185493
R1997 X1.n171 X1.n170 0.00184889
R1998 X1.n180 X1.n95 0.00184889
R1999 X1.n798 X1.n464 0.00184889
R2000 X1.n1018 X1.n365 0.00184889
R2001 X1.n1097 X1.n1095 0.00184889
R2002 X1.n1193 X1.n1192 0.00184889
R2003 X1.n1202 X1.n1201 0.00184889
R2004 X1.n1293 X1.n1292 0.00184889
R2005 X1.n554 X1.n553 0.00184889
R2006 X1.n746 X1.n495 0.00184889
R2007 X1.n736 X1.n625 0.00184889
R2008 X1.n669 X1.n667 0.00184889
R2009 X1.n997 X1.n373 0.00183571
R2010 X1.n1049 X1.n1044 0.00182678
R2011 X1.n859 X1.n437 0.00180952
R2012 X1.n143 X1.n48 0.0017973
R2013 X1.n207 X1.n64 0.0017973
R2014 X1.n855 X1.n439 0.0017973
R2015 X1.n1001 X1.n371 0.0017973
R2016 X1.n557 X1.n526 0.0017897
R2017 X1.n733 X1.n732 0.0017897
R2018 X1.n887 X1.n422 0.00178256
R2019 X1.n894 X1.n893 0.00178256
R2020 X1.n972 X1.n971 0.00178256
R2021 X1.n960 X1.n392 0.00176044
R2022 X1.n677 X1.n676 0.00175714
R2023 X1.n861 X1.n860 0.00173095
R2024 X1.n996 X1.n995 0.00173095
R2025 X1.n807 X1.n806 0.00171622
R2026 X1.n620 X1.n503 0.00171347
R2027 X1.n1343 X1.n1342 0.0016941
R2028 X1.n244 X1.n82 0.0016941
R2029 X1.n829 X1.n450 0.0016941
R2030 X1.n363 X1.n360 0.0016941
R2031 X1.n1058 X1.n1039 0.0016941
R2032 X1.n1031 X1.n1030 0.00165238
R2033 X1.n917 X1.n916 0.00162776
R2034 X1.n924 X1.n923 0.00162776
R2035 X1.n998 X1.n374 0.00162776
R2036 X1.n1092 X1.n1091 0.00162776
R2037 X1.n826 X1.n825 0.00162619
R2038 X1.n858 X1.n438 0.00160565
R2039 X1.n1116 X1.n1115 0.00158354
R2040 X1.n289 X1.n288 0.00158354
R2041 X1.n567 X1.n566 0.00158354
R2042 X1.n728 X1.n628 0.00158354
R2043 X1.n162 X1.n99 0.00156143
R2044 X1.n187 X1.n94 0.00156143
R2045 X1.n797 X1.n796 0.00156143
R2046 X1.n1048 X1.n1047 0.00156143
R2047 X1.n1174 X1.n1173 0.00156143
R2048 X1.n1279 X1.n1278 0.00156143
R2049 X1.n622 X1.n501 0.00156143
R2050 X1.n675 X1.n662 0.00156143
R2051 X1.n896 X1.n416 0.00154762
R2052 X1.n957 X1.n393 0.00154762
R2053 X1.n862 X1.n436 0.00153931
R2054 X1.n994 X1.n376 0.00153931
R2055 X1.n897 X1.n417 0.00149509
R2056 X1.n659 X1.n658 0.00149509
R2057 X1.n956 X1.n955 0.00147297
R2058 X1.n1029 X1.n357 0.00147297
R2059 X1.n794 X1.n466 0.00146905
R2060 X1.n1046 X1.n1045 0.00146905
R2061 X1.n824 X1.n452 0.00145086
R2062 X1.n125 X1.n108 0.00140663
R2063 X1.n226 X1.n85 0.00140663
R2064 X1.n830 X1.n452 0.00140663
R2065 X1.n1029 X1.n1028 0.00140663
R2066 X1.n922 X1.n921 0.00139048
R2067 X1.n898 X1.n897 0.00138452
R2068 X1.n956 X1.n394 0.00138452
R2069 X1.n535 X1.n534 0.00136429
R2070 X1.n903 X1.n902 0.00136429
R2071 X1.n914 X1.n409 0.00136429
R2072 X1.n857 X1.n436 0.00134029
R2073 X1.n999 X1.n376 0.00134029
R2074 X1.n944 X1.n397 0.00133809
R2075 X1.n1080 X1.n344 0.00133809
R2076 X1.n796 X1.n795 0.00131818
R2077 X1.n1047 X1.n347 0.00131818
R2078 X1.n622 X1.n621 0.00131818
R2079 X1.n1138 X1.n1137 0.00129607
R2080 X1.n1162 X1.n1161 0.00129607
R2081 X1.n1221 X1.n1220 0.00129607
R2082 X1.n1254 X1.n1251 0.00129607
R2083 X1.n809 X1.n808 0.00128571
R2084 X1.n1057 X1.n1038 0.00128571
R2085 X1.n147 X1.n146 0.00125184
R2086 X1.n204 X1.n203 0.00125184
R2087 X1.n858 X1.n857 0.00125184
R2088 X1.n923 X1.n400 0.00125184
R2089 X1.n999 X1.n998 0.00125184
R2090 X1.n537 X1.n469 0.00122973
R2091 X1.n415 X1.n412 0.00122973
R2092 X1.n916 X1.n915 0.00122973
R2093 X1.n946 X1.n945 0.00120762
R2094 X1.n1082 X1.n1081 0.00120762
R2095 X1.n868 X1.n421 0.00120714
R2096 X1.n970 X1.n969 0.00120714
R2097 X1.n830 X1.n829 0.0011855
R2098 X1.n1028 X1.n360 0.0011855
R2099 X1.n807 X1.n460 0.00116339
R2100 X1.n1059 X1.n1058 0.00116339
R2101 X1.n1126 X1.n328 0.00114865
R2102 X1.n1213 X1.n1212 0.00114865
R2103 X1.n562 X1.n479 0.00114865
R2104 X1.n725 X1.n630 0.00114865
R2105 X1.n1013 X1.n364 0.00112857
R2106 X1.n955 X1.n392 0.00111916
R2107 X1.n837 X1.n445 0.00110238
R2108 X1.n142 X1.n141 0.00109705
R2109 X1.n209 X1.n208 0.00109705
R2110 X1.n869 X1.n422 0.00109705
R2111 X1.n894 X1.n417 0.00109705
R2112 X1.n971 X1.n390 0.00109705
R2113 X1.n680 X1.n658 0.00109705
R2114 X1.n1142 X1.n309 0.00105283
R2115 X1.n1256 X1.n1249 0.00105283
R2116 X1.n247 X1.n79 0.00105283
R2117 X1.n168 X1.n55 0.00104054
R2118 X1.n931 X1.n405 0.00104054
R2119 X1.n798 X1.n797 0.00103071
R2120 X1.n368 X1.n365 0.00103071
R2121 X1.n1049 X1.n1048 0.00103071
R2122 X1.n1088 X1.n341 0.00103071
R2123 X1.n322 X1.n316 0.00103071
R2124 X1.n1239 X1.n1238 0.00103071
R2125 X1.n542 X1.n530 0.00103071
R2126 X1.n555 X1.n554 0.00103071
R2127 X1.n626 X1.n625 0.00103071
R2128 X1.n838 X1.n446 0.0010086
R2129 X1.n918 X1.n917 0.000964373
R2130 X1.n925 X1.n924 0.000964373
R2131 X1.n1091 X1.n342 0.000964373
R2132 X1.n549 X1.n547 0.000964373
R2133 X1.n668 X1.n31 0.000964373
R2134 X1.n130 X1.n129 0.00094226
R2135 X1.n219 X1.n86 0.00094226
R2136 X1.n1122 X1.n329 0.000932432
R2137 X1.n1227 X1.n1226 0.000932432
R2138 X1.n575 X1.n480 0.000932432
R2139 X1.n714 X1.n12 0.000932432
R2140 X1.n543 X1.n529 0.000898034
R2141 X1.n1055 X1.n1039 0.000898034
R2142 X1.n806 X1.n462 0.000875921
R2143 X1.n1103 X1.n340 0.000853808
R2144 X1.n684 X1.n654 0.000831695
R2145 X1.n657 X1.n656 0.000814286
R2146 X1.n888 X1.n887 0.000809582
R2147 X1.n972 X1.n389 0.000809582
R2148 X1.n155 X1.n100 0.000787469
R2149 X1.n192 X1.n191 0.000787469
R2150 X1.n579 X1.n578 0.000787469
R2151 X1.n718 X1.n717 0.000787469
R2152 X1.n1119 X1.n330 0.000765356
R2153 X1.n1177 X1.n305 0.000765356
R2154 X1.n1215 X1.n1214 0.000765356
R2155 X1.n1274 X1.n1273 0.000765356
R2156 X1.n681 X1.n655 0.000765356
R2157 X1.n1019 X1.n1018 0.000743243
R2158 X1.n839 X1.n448 0.00072113
R2159 X1.n116 X1.n112 0.000716216
R2160 X1.n234 X1.n70 0.000716216
R2161 X1.n805 X1.n459 0.000716216
R2162 X1.n1042 X1.n1041 0.000716216
R2163 X1.n850 X1.n849 0.000676904
R2164 X1.n114 X1.n113 0.000654791
R2165 X1.n237 X1.n236 0.000654791
R2166 X1.n1007 X1.n1006 0.000654791
R2167 X1.n987 X1.n378 0.000588452
R2168 X1.n876 X1.n433 0.000566339
R2169 X1.n1347 X1.n30 0.000522113
R2170 X1.n820 X1.n819 0.000522113
R2171 X2.n3 X2.n0 15.1893
R2172 X2.n2 X2.n1 15.0005
R2173 X2.n4 X2.n3 9.50738
R2174 X2.n1378 X2.n4 9.08058
R2175 X2.n1378 X2 2.85925
R2176 X2.n605 X2.n51 2.2505
R2177 X2.n1326 X2.n49 2.2505
R2178 X2.n624 X2.n46 2.2505
R2179 X2.n1332 X2.n44 2.2505
R2180 X2.n642 X2.n41 2.2505
R2181 X2.n1338 X2.n39 2.2505
R2182 X2.n576 X2.n36 2.2505
R2183 X2.n1343 X2.n35 2.2505
R2184 X2.n1345 X2.n33 2.2505
R2185 X2.n1349 X2.n30 2.2505
R2186 X2.n1351 X2.n28 2.2505
R2187 X2.n1355 X2.n25 2.2505
R2188 X2.n1357 X2.n23 2.2505
R2189 X2.n1361 X2.n20 2.2505
R2190 X2.n1363 X2.n18 2.2505
R2191 X2.n1323 X2.n51 2.2505
R2192 X2.n1326 X2.n47 2.2505
R2193 X2.n1329 X2.n46 2.2505
R2194 X2.n1332 X2.n42 2.2505
R2195 X2.n1335 X2.n41 2.2505
R2196 X2.n1338 X2.n37 2.2505
R2197 X2.n1341 X2.n36 2.2505
R2198 X2.n1343 X2.n1342 2.2505
R2199 X2.n1346 X2.n1345 2.2505
R2200 X2.n1349 X2.n1348 2.2505
R2201 X2.n1352 X2.n1351 2.2505
R2202 X2.n1355 X2.n1354 2.2505
R2203 X2.n1358 X2.n1357 2.2505
R2204 X2.n1361 X2.n1360 2.2505
R2205 X2.n1364 X2.n1363 2.2505
R2206 X2.n282 X2.n281 2.2505
R2207 X2.n283 X2.n270 2.2505
R2208 X2.n805 X2.n262 2.2505
R2209 X2.n801 X2.n254 2.2505
R2210 X2.n903 X2.n902 2.2505
R2211 X2.n909 X2.n908 2.2505
R2212 X2.n931 X2.n215 2.2505
R2213 X2.n213 X2.n212 2.2505
R2214 X2.n961 X2.n960 2.2505
R2215 X2.n999 X2.n998 2.2505
R2216 X2.n1009 X2.n1008 2.2505
R2217 X2.n1004 X2.n177 2.2505
R2218 X2.n1050 X2.n162 2.2505
R2219 X2.n1065 X2.n160 2.2505
R2220 X2.n1097 X2.n148 2.2505
R2221 X2.n799 X2.n282 2.2505
R2222 X2.n808 X2.n283 2.2505
R2223 X2.n805 X2.n800 2.2505
R2224 X2.n802 X2.n801 2.2505
R2225 X2.n904 X2.n903 2.2505
R2226 X2.n908 X2.n907 2.2505
R2227 X2.n215 X2.n214 2.2505
R2228 X2.n958 X2.n213 2.2505
R2229 X2.n960 X2.n959 2.2505
R2230 X2.n1000 X2.n999 2.2505
R2231 X2.n1008 X2.n1007 2.2505
R2232 X2.n1005 X2.n1004 2.2505
R2233 X2.n162 X2.n161 2.2505
R2234 X2.n1093 X2.n160 2.2505
R2235 X2.n148 X2.n147 2.2505
R2236 X2.n53 X2.n52 2.2505
R2237 X2.n1311 X2.n1310 2.2505
R2238 X2.n1309 X2.n63 2.2505
R2239 X2.n1308 X2.n1307 2.2505
R2240 X2.n65 X2.n64 2.2505
R2241 X2.n1287 X2.n1286 2.2505
R2242 X2.n1285 X2.n72 2.2505
R2243 X2.n1284 X2.n1283 2.2505
R2244 X2.n74 X2.n73 2.2505
R2245 X2.n1257 X2.n1256 2.2505
R2246 X2.n1258 X2.n1255 2.2505
R2247 X2.n1254 X2.n83 2.2505
R2248 X2.n1253 X2.n1252 2.2505
R2249 X2.n85 X2.n84 2.2505
R2250 X2.n1233 X2.n1232 2.2505
R2251 X2.n1231 X2.n93 2.2505
R2252 X2.n1230 X2.n1229 2.2505
R2253 X2.n95 X2.n94 2.2505
R2254 X2.n1210 X2.n1209 2.2505
R2255 X2.n1211 X2.n1208 2.2505
R2256 X2.n1207 X2.n110 2.2505
R2257 X2.n1206 X2.n1205 2.2505
R2258 X2.n112 X2.n111 2.2505
R2259 X2.n1179 X2.n1178 2.2505
R2260 X2.n1180 X2.n1177 2.2505
R2261 X2.n1176 X2.n122 2.2505
R2262 X2.n1175 X2.n1174 2.2505
R2263 X2.n124 X2.n123 2.2505
R2264 X2.n1155 X2.n1154 2.2505
R2265 X2.n1153 X2.n136 2.2505
R2266 X2.n1152 X2.n1151 2.2505
R2267 X2.n138 X2.n137 2.2505
R2268 X2.n1133 X2.n1132 2.2505
R2269 X2.n1131 X2.n146 2.2505
R2270 X2.n1117 X2.n146 2.2505
R2271 X2.n1134 X2.n1133 2.2505
R2272 X2.n1137 X2.n138 2.2505
R2273 X2.n1151 X2.n1150 2.2505
R2274 X2.n140 X2.n136 2.2505
R2275 X2.n1156 X2.n1155 2.2505
R2276 X2.n1159 X2.n124 2.2505
R2277 X2.n1174 X2.n1173 2.2505
R2278 X2.n128 X2.n122 2.2505
R2279 X2.n1181 X2.n1180 2.2505
R2280 X2.n1179 X2.n119 2.2505
R2281 X2.n1189 X2.n112 2.2505
R2282 X2.n1205 X2.n1204 2.2505
R2283 X2.n1194 X2.n110 2.2505
R2284 X2.n1212 X2.n1211 2.2505
R2285 X2.n1210 X2.n107 2.2505
R2286 X2.n1220 X2.n95 2.2505
R2287 X2.n1229 X2.n1228 2.2505
R2288 X2.n101 X2.n93 2.2505
R2289 X2.n1234 X2.n1233 2.2505
R2290 X2.n1236 X2.n85 2.2505
R2291 X2.n1252 X2.n1251 2.2505
R2292 X2.n1241 X2.n83 2.2505
R2293 X2.n1259 X2.n1258 2.2505
R2294 X2.n1257 X2.n80 2.2505
R2295 X2.n1267 X2.n74 2.2505
R2296 X2.n1283 X2.n1282 2.2505
R2297 X2.n1276 X2.n72 2.2505
R2298 X2.n1288 X2.n1287 2.2505
R2299 X2.n1291 X2.n65 2.2505
R2300 X2.n1307 X2.n1306 2.2505
R2301 X2.n1299 X2.n63 2.2505
R2302 X2.n1312 X2.n1311 2.2505
R2303 X2.n55 X2.n53 2.2505
R2304 X2.n796 X2.n286 2.2505
R2305 X2.n795 X2.n287 2.2505
R2306 X2.n409 X2.n288 2.2505
R2307 X2.n791 X2.n290 2.2505
R2308 X2.n790 X2.n291 2.2505
R2309 X2.n789 X2.n292 2.2505
R2310 X2.n361 X2.n293 2.2505
R2311 X2.n785 X2.n295 2.2505
R2312 X2.n784 X2.n296 2.2505
R2313 X2.n783 X2.n297 2.2505
R2314 X2.n356 X2.n298 2.2505
R2315 X2.n779 X2.n300 2.2505
R2316 X2.n778 X2.n301 2.2505
R2317 X2.n777 X2.n302 2.2505
R2318 X2.n350 X2.n303 2.2505
R2319 X2.n773 X2.n305 2.2505
R2320 X2.n772 X2.n306 2.2505
R2321 X2.n771 X2.n307 2.2505
R2322 X2.n494 X2.n308 2.2505
R2323 X2.n767 X2.n310 2.2505
R2324 X2.n766 X2.n311 2.2505
R2325 X2.n765 X2.n312 2.2505
R2326 X2.n508 X2.n313 2.2505
R2327 X2.n761 X2.n315 2.2505
R2328 X2.n760 X2.n316 2.2505
R2329 X2.n759 X2.n757 2.2505
R2330 X2.n517 X2.n7 2.2505
R2331 X2.n1375 X2.n8 2.2505
R2332 X2.n1374 X2.n9 2.2505
R2333 X2.n1373 X2.n10 2.2505
R2334 X2.n530 X2.n11 2.2505
R2335 X2.n1369 X2.n13 2.2505
R2336 X2.n1368 X2.n14 2.2505
R2337 X2.n1367 X2.n15 2.2505
R2338 X2.n1367 X2.n1366 2.2505
R2339 X2.n1368 X2.n12 2.2505
R2340 X2.n1370 X2.n1369 2.2505
R2341 X2.n1371 X2.n11 2.2505
R2342 X2.n1373 X2.n1372 2.2505
R2343 X2.n1374 X2.n6 2.2505
R2344 X2.n1376 X2.n1375 2.2505
R2345 X2.n7 X2.n5 2.2505
R2346 X2.n759 X2.n758 2.2505
R2347 X2.n760 X2.n314 2.2505
R2348 X2.n762 X2.n761 2.2505
R2349 X2.n763 X2.n313 2.2505
R2350 X2.n765 X2.n764 2.2505
R2351 X2.n766 X2.n309 2.2505
R2352 X2.n768 X2.n767 2.2505
R2353 X2.n769 X2.n308 2.2505
R2354 X2.n771 X2.n770 2.2505
R2355 X2.n772 X2.n304 2.2505
R2356 X2.n774 X2.n773 2.2505
R2357 X2.n775 X2.n303 2.2505
R2358 X2.n777 X2.n776 2.2505
R2359 X2.n778 X2.n299 2.2505
R2360 X2.n780 X2.n779 2.2505
R2361 X2.n781 X2.n298 2.2505
R2362 X2.n783 X2.n782 2.2505
R2363 X2.n784 X2.n294 2.2505
R2364 X2.n786 X2.n785 2.2505
R2365 X2.n787 X2.n293 2.2505
R2366 X2.n789 X2.n788 2.2505
R2367 X2.n790 X2.n289 2.2505
R2368 X2.n792 X2.n791 2.2505
R2369 X2.n793 X2.n288 2.2505
R2370 X2.n795 X2.n794 2.2505
R2371 X2.n796 X2.n284 2.2505
R2372 X2.n56 X2.n54 2.2005
R2373 X2.n725 X2.n724 2.2005
R2374 X2.n723 X2.n722 2.2005
R2375 X2.n721 X2.n720 2.2005
R2376 X2.n719 X2.n718 2.2005
R2377 X2.n717 X2.n548 2.2005
R2378 X2.n716 X2.n715 2.2005
R2379 X2.n714 X2.n713 2.2005
R2380 X2.n712 X2.n711 2.2005
R2381 X2.n710 X2.n709 2.2005
R2382 X2.n708 X2.n707 2.2005
R2383 X2.n706 X2.n705 2.2005
R2384 X2.n704 X2.n703 2.2005
R2385 X2.n559 X2.n553 2.2005
R2386 X2.n561 X2.n560 2.2005
R2387 X2.n698 X2.n697 2.2005
R2388 X2.n696 X2.n562 2.2005
R2389 X2.n694 X2.n693 2.2005
R2390 X2.n692 X2.n563 2.2005
R2391 X2.n691 X2.n690 2.2005
R2392 X2.n567 X2.n565 2.2005
R2393 X2.n569 X2.n568 2.2005
R2394 X2.n685 X2.n684 2.2005
R2395 X2.n683 X2.n682 2.2005
R2396 X2.n680 X2.n679 2.2005
R2397 X2.n678 X2.n570 2.2005
R2398 X2.n676 X2.n675 2.2005
R2399 X2.n572 X2.n571 2.2005
R2400 X2.n667 X2.n574 2.2005
R2401 X2.n670 X2.n669 2.2005
R2402 X2.n668 X2.n666 2.2005
R2403 X2.n665 X2.n664 2.2005
R2404 X2.n663 X2.n662 2.2005
R2405 X2.n661 X2.n660 2.2005
R2406 X2.n659 X2.n658 2.2005
R2407 X2.n657 X2.n656 2.2005
R2408 X2.n655 X2.n654 2.2005
R2409 X2.n653 X2.n652 2.2005
R2410 X2.n651 X2.n650 2.2005
R2411 X2.n582 X2.n578 2.2005
R2412 X2.n584 X2.n583 2.2005
R2413 X2.n645 X2.n644 2.2005
R2414 X2.n643 X2.n585 2.2005
R2415 X2.n641 X2.n640 2.2005
R2416 X2.n639 X2.n586 2.2005
R2417 X2.n638 X2.n637 2.2005
R2418 X2.n590 X2.n588 2.2005
R2419 X2.n592 X2.n591 2.2005
R2420 X2.n632 X2.n631 2.2005
R2421 X2.n630 X2.n629 2.2005
R2422 X2.n627 X2.n626 2.2005
R2423 X2.n625 X2.n593 2.2005
R2424 X2.n623 X2.n622 2.2005
R2425 X2.n595 X2.n594 2.2005
R2426 X2.n615 X2.n597 2.2005
R2427 X2.n617 X2.n616 2.2005
R2428 X2.n614 X2.n613 2.2005
R2429 X2.n612 X2.n611 2.2005
R2430 X2.n610 X2.n599 2.2005
R2431 X2.n609 X2.n608 2.2005
R2432 X2.n607 X2.n606 2.2005
R2433 X2.n1107 X2.n149 2.2005
R2434 X2.n1098 X2.n156 2.2005
R2435 X2.n1100 X2.n1099 2.2005
R2436 X2.n1072 X2.n159 2.2005
R2437 X2.n1077 X2.n1067 2.2005
R2438 X2.n1066 X2.n1063 2.2005
R2439 X2.n1084 X2.n164 2.2005
R2440 X2.n1089 X2.n1088 2.2005
R2441 X2.n1059 X2.n163 2.2005
R2442 X2.n1057 X2.n169 2.2005
R2443 X2.n1052 X2.n1051 2.2005
R2444 X2.n1049 X2.n1048 2.2005
R2445 X2.n1042 X2.n1041 2.2005
R2446 X2.n1040 X2.n1039 2.2005
R2447 X2.n1034 X2.n1033 2.2005
R2448 X2.n1032 X2.n1031 2.2005
R2449 X2.n1026 X2.n1025 2.2005
R2450 X2.n1024 X2.n1023 2.2005
R2451 X2.n1017 X2.n186 2.2005
R2452 X2.n1011 X2.n1010 2.2005
R2453 X2.n192 X2.n191 2.2005
R2454 X2.n991 X2.n199 2.2005
R2455 X2.n997 X2.n996 2.2005
R2456 X2.n985 X2.n197 2.2005
R2457 X2.n979 X2.n978 2.2005
R2458 X2.n976 X2.n975 2.2005
R2459 X2.n971 X2.n206 2.2005
R2460 X2.n962 X2.n209 2.2005
R2461 X2.n964 X2.n963 2.2005
R2462 X2.n948 X2.n217 2.2005
R2463 X2.n954 X2.n953 2.2005
R2464 X2.n941 X2.n216 2.2005
R2465 X2.n932 X2.n221 2.2005
R2466 X2.n934 X2.n933 2.2005
R2467 X2.n930 X2.n929 2.2005
R2468 X2.n923 X2.n224 2.2005
R2469 X2.n236 X2.n228 2.2005
R2470 X2.n916 X2.n231 2.2005
R2471 X2.n911 X2.n910 2.2005
R2472 X2.n894 X2.n234 2.2005
R2473 X2.n245 X2.n243 2.2005
R2474 X2.n901 X2.n900 2.2005
R2475 X2.n887 X2.n241 2.2005
R2476 X2.n881 X2.n880 2.2005
R2477 X2.n879 X2.n878 2.2005
R2478 X2.n873 X2.n872 2.2005
R2479 X2.n871 X2.n870 2.2005
R2480 X2.n866 X2.n865 2.2005
R2481 X2.n864 X2.n863 2.2005
R2482 X2.n857 X2.n856 2.2005
R2483 X2.n855 X2.n854 2.2005
R2484 X2.n847 X2.n846 2.2005
R2485 X2.n845 X2.n844 2.2005
R2486 X2.n838 X2.n837 2.2005
R2487 X2.n836 X2.n835 2.2005
R2488 X2.n830 X2.n829 2.2005
R2489 X2.n828 X2.n827 2.2005
R2490 X2.n821 X2.n274 2.2005
R2491 X2.n812 X2.n278 2.2005
R2492 X2.n814 X2.n813 2.2005
R2493 X2.n383 X2.n381 2.2005
R2494 X2.n1115 X2.n150 2.2005
R2495 X2.n1119 X2.n1118 2.2005
R2496 X2.n1120 X2.n145 2.2005
R2497 X2.n1135 X2.n143 2.2005
R2498 X2.n1139 X2.n1138 2.2005
R2499 X2.n1136 X2.n144 2.2005
R2500 X2.n141 X2.n139 2.2005
R2501 X2.n1149 X2.n1148 2.2005
R2502 X2.n1147 X2.n1146 2.2005
R2503 X2.n1144 X2.n135 2.2005
R2504 X2.n1157 X2.n132 2.2005
R2505 X2.n1161 X2.n1160 2.2005
R2506 X2.n1158 X2.n134 2.2005
R2507 X2.n133 X2.n125 2.2005
R2508 X2.n1172 X2.n1171 2.2005
R2509 X2.n1170 X2.n126 2.2005
R2510 X2.n130 X2.n129 2.2005
R2511 X2.n1165 X2.n121 2.2005
R2512 X2.n1182 X2.n120 2.2005
R2513 X2.n1184 X2.n1183 2.2005
R2514 X2.n1187 X2.n1186 2.2005
R2515 X2.n1188 X2.n118 2.2005
R2516 X2.n1191 X2.n1190 2.2005
R2517 X2.n115 X2.n113 2.2005
R2518 X2.n1203 X2.n1202 2.2005
R2519 X2.n116 X2.n114 2.2005
R2520 X2.n1196 X2.n1195 2.2005
R2521 X2.n1197 X2.n109 2.2005
R2522 X2.n1213 X2.n108 2.2005
R2523 X2.n1215 X2.n1214 2.2005
R2524 X2.n1218 X2.n1217 2.2005
R2525 X2.n1219 X2.n106 2.2005
R2526 X2.n1222 X2.n1221 2.2005
R2527 X2.n98 X2.n96 2.2005
R2528 X2.n1227 X2.n1226 2.2005
R2529 X2.n104 X2.n97 2.2005
R2530 X2.n103 X2.n102 2.2005
R2531 X2.n99 X2.n92 2.2005
R2532 X2.n1235 X2.n91 2.2005
R2533 X2.n1238 X2.n1237 2.2005
R2534 X2.n88 X2.n86 2.2005
R2535 X2.n1250 X2.n1249 2.2005
R2536 X2.n89 X2.n87 2.2005
R2537 X2.n1243 X2.n1242 2.2005
R2538 X2.n1244 X2.n82 2.2005
R2539 X2.n1260 X2.n81 2.2005
R2540 X2.n1262 X2.n1261 2.2005
R2541 X2.n1265 X2.n1264 2.2005
R2542 X2.n1266 X2.n79 2.2005
R2543 X2.n1269 X2.n1268 2.2005
R2544 X2.n77 X2.n75 2.2005
R2545 X2.n1281 X2.n1280 2.2005
R2546 X2.n1279 X2.n76 2.2005
R2547 X2.n1278 X2.n1277 2.2005
R2548 X2.n1274 X2.n71 2.2005
R2549 X2.n1289 X2.n70 2.2005
R2550 X2.n1293 X2.n1292 2.2005
R2551 X2.n1290 X2.n68 2.2005
R2552 X2.n1298 X2.n66 2.2005
R2553 X2.n1305 X2.n1304 2.2005
R2554 X2.n1303 X2.n67 2.2005
R2555 X2.n1301 X2.n1300 2.2005
R2556 X2.n62 X2.n61 2.2005
R2557 X2.n1315 X2.n1314 2.2005
R2558 X2.n1313 X2.n57 2.2005
R2559 X2.n394 X2.n393 2.2005
R2560 X2.n398 X2.n397 2.2005
R2561 X2.n396 X2.n371 2.2005
R2562 X2.n405 X2.n403 2.2005
R2563 X2.n411 X2.n410 2.2005
R2564 X2.n408 X2.n404 2.2005
R2565 X2.n407 X2.n406 2.2005
R2566 X2.n368 X2.n367 2.2005
R2567 X2.n420 X2.n415 2.2005
R2568 X2.n422 X2.n421 2.2005
R2569 X2.n418 X2.n417 2.2005
R2570 X2.n416 X2.n362 2.2005
R2571 X2.n429 X2.n428 2.2005
R2572 X2.n431 X2.n430 2.2005
R2573 X2.n434 X2.n433 2.2005
R2574 X2.n436 X2.n435 2.2005
R2575 X2.n439 X2.n438 2.2005
R2576 X2.n437 X2.n358 2.2005
R2577 X2.n445 X2.n444 2.2005
R2578 X2.n447 X2.n446 2.2005
R2579 X2.n450 X2.n449 2.2005
R2580 X2.n452 X2.n451 2.2005
R2581 X2.n457 X2.n453 2.2005
R2582 X2.n459 X2.n458 2.2005
R2583 X2.n456 X2.n455 2.2005
R2584 X2.n454 X2.n352 2.2005
R2585 X2.n465 X2.n464 2.2005
R2586 X2.n467 X2.n466 2.2005
R2587 X2.n472 X2.n471 2.2005
R2588 X2.n474 X2.n473 2.2005
R2589 X2.n477 X2.n476 2.2005
R2590 X2.n475 X2.n347 2.2005
R2591 X2.n483 X2.n482 2.2005
R2592 X2.n485 X2.n484 2.2005
R2593 X2.n487 X2.n345 2.2005
R2594 X2.n493 X2.n492 2.2005
R2595 X2.n495 X2.n340 2.2005
R2596 X2.n497 X2.n496 2.2005
R2597 X2.n344 X2.n343 2.2005
R2598 X2.n342 X2.n341 2.2005
R2599 X2.n337 X2.n336 2.2005
R2600 X2.n503 X2.n501 2.2005
R2601 X2.n510 X2.n509 2.2005
R2602 X2.n507 X2.n506 2.2005
R2603 X2.n505 X2.n504 2.2005
R2604 X2.n331 X2.n330 2.2005
R2605 X2.n329 X2.n328 2.2005
R2606 X2.n325 X2.n324 2.2005
R2607 X2.n323 X2.n317 2.2005
R2608 X2.n756 X2.n755 2.2005
R2609 X2.n754 X2.n318 2.2005
R2610 X2.n518 X2.n320 2.2005
R2611 X2.n520 X2.n519 2.2005
R2612 X2.n525 X2.n524 2.2005
R2613 X2.n527 X2.n526 2.2005
R2614 X2.n746 X2.n528 2.2005
R2615 X2.n748 X2.n747 2.2005
R2616 X2.n745 X2.n744 2.2005
R2617 X2.n743 X2.n742 2.2005
R2618 X2.n536 X2.n534 2.2005
R2619 X2.n538 X2.n537 2.2005
R2620 X2.n735 X2.n734 2.2005
R2621 X2.n733 X2.n732 2.2005
R2622 X2.n541 X2.n540 2.2005
R2623 X2.n543 X2.n542 2.2005
R2624 X2.n1325 X2.n50 1.8005
R2625 X2.n1327 X2.n48 1.8005
R2626 X2.n1331 X2.n45 1.8005
R2627 X2.n1333 X2.n43 1.8005
R2628 X2.n1337 X2.n40 1.8005
R2629 X2.n1339 X2.n38 1.8005
R2630 X2.n1344 X2.n34 1.8005
R2631 X2.n677 X2.n31 1.8005
R2632 X2.n1350 X2.n29 1.8005
R2633 X2.n695 X2.n26 1.8005
R2634 X2.n1356 X2.n24 1.8005
R2635 X2.n551 X2.n21 1.8005
R2636 X2.n1362 X2.n19 1.8005
R2637 X2.n1325 X2.n1324 1.8005
R2638 X2.n1328 X2.n1327 1.8005
R2639 X2.n1331 X2.n1330 1.8005
R2640 X2.n1334 X2.n1333 1.8005
R2641 X2.n1337 X2.n1336 1.8005
R2642 X2.n1340 X2.n1339 1.8005
R2643 X2.n1344 X2.n32 1.8005
R2644 X2.n1347 X2.n31 1.8005
R2645 X2.n1350 X2.n27 1.8005
R2646 X2.n1353 X2.n26 1.8005
R2647 X2.n1356 X2.n22 1.8005
R2648 X2.n1359 X2.n21 1.8005
R2649 X2.n1362 X2.n17 1.8005
R2650 X2.n811 X2.n810 1.8005
R2651 X2.n806 X2.n266 1.8005
R2652 X2.n804 X2.n258 1.8005
R2653 X2.n250 X2.n240 1.8005
R2654 X2.n242 X2.n235 1.8005
R2655 X2.n238 X2.n237 1.8005
R2656 X2.n956 X2.n955 1.8005
R2657 X2.n977 X2.n196 1.8005
R2658 X2.n198 X2.n193 1.8005
R2659 X2.n194 X2.n182 1.8005
R2660 X2.n1003 X2.n172 1.8005
R2661 X2.n1091 X2.n1090 1.8005
R2662 X2.n1096 X2.n1095 1.8005
R2663 X2.n810 X2.n809 1.8005
R2664 X2.n807 X2.n806 1.8005
R2665 X2.n804 X2.n803 1.8005
R2666 X2.n240 X2.n239 1.8005
R2667 X2.n905 X2.n235 1.8005
R2668 X2.n906 X2.n238 1.8005
R2669 X2.n957 X2.n956 1.8005
R2670 X2.n196 X2.n195 1.8005
R2671 X2.n1001 X2.n193 1.8005
R2672 X2.n1006 X2.n194 1.8005
R2673 X2.n1003 X2.n1002 1.8005
R2674 X2.n1092 X2.n1091 1.8005
R2675 X2.n1095 X2.n1094 1.8005
R2676 X2.n1322 X2.n1321 1.8005
R2677 X2.n1321 X2.n1320 1.8005
R2678 X2.n726 X2.n16 1.8005
R2679 X2.n1365 X2.n16 1.8005
R2680 X2.n1130 X2.n1129 1.5005
R2681 X2.n1129 X2.n1128 1.5005
R2682 X2.n797 X2.n285 1.5005
R2683 X2.n798 X2.n797 1.5005
R2684 X2.n1124 X2.n1116 1.1125
R2685 X2.n739 X2.n535 1.10836
R2686 X2.n741 X2.n740 1.10443
R2687 X2.n729 X2.n544 1.10381
R2688 X2.n1125 X2.n153 1.10372
R2689 X2.n529 X2.n523 1.10339
R2690 X2.n735 X2.n539 1.10272
R2691 X2.n738 X2.n538 1.10272
R2692 X2.n742 X2.n533 1.10272
R2693 X2.n1123 X2.n1119 1.10263
R2694 X2.n1120 X2.n142 1.10263
R2695 X2.n604 X2.n603 1.1005
R2696 X2.n554 X2.n547 1.1005
R2697 X2.n555 X2.n549 1.1005
R2698 X2.n556 X2.n550 1.1005
R2699 X2.n557 X2.n552 1.1005
R2700 X2.n702 X2.n701 1.1005
R2701 X2.n700 X2.n699 1.1005
R2702 X2.n564 X2.n558 1.1005
R2703 X2.n689 X2.n688 1.1005
R2704 X2.n687 X2.n686 1.1005
R2705 X2.n681 X2.n566 1.1005
R2706 X2.n674 X2.n673 1.1005
R2707 X2.n672 X2.n671 1.1005
R2708 X2.n665 X2.n573 1.1005
R2709 X2.n579 X2.n575 1.1005
R2710 X2.n580 X2.n577 1.1005
R2711 X2.n649 X2.n648 1.1005
R2712 X2.n647 X2.n646 1.1005
R2713 X2.n587 X2.n581 1.1005
R2714 X2.n636 X2.n635 1.1005
R2715 X2.n634 X2.n633 1.1005
R2716 X2.n628 X2.n589 1.1005
R2717 X2.n621 X2.n620 1.1005
R2718 X2.n619 X2.n618 1.1005
R2719 X2.n598 X2.n596 1.1005
R2720 X2.n546 X2.n545 1.1005
R2721 X2.n600 X2.n58 1.1005
R2722 X2.n601 X2.n59 1.1005
R2723 X2.n602 X2.n601 1.1005
R2724 X2.n1319 X2.n1318 1.1005
R2725 X2.n1317 X2.n1316 1.1005
R2726 X2.n1302 X2.n60 1.1005
R2727 X2.n1297 X2.n1296 1.1005
R2728 X2.n1295 X2.n1294 1.1005
R2729 X2.n1275 X2.n69 1.1005
R2730 X2.n1273 X2.n1272 1.1005
R2731 X2.n1271 X2.n1270 1.1005
R2732 X2.n1263 X2.n78 1.1005
R2733 X2.n1246 X2.n1245 1.1005
R2734 X2.n1248 X2.n1247 1.1005
R2735 X2.n1240 X2.n1239 1.1005
R2736 X2.n100 X2.n90 1.1005
R2737 X2.n1225 X2.n1224 1.1005
R2738 X2.n1223 X2.n1222 1.1005
R2739 X2.n1216 X2.n105 1.1005
R2740 X2.n1199 X2.n1198 1.1005
R2741 X2.n1201 X2.n1200 1.1005
R2742 X2.n1193 X2.n1192 1.1005
R2743 X2.n1185 X2.n117 1.1005
R2744 X2.n1167 X2.n1166 1.1005
R2745 X2.n1169 X2.n1168 1.1005
R2746 X2.n1164 X2.n127 1.1005
R2747 X2.n1163 X2.n1162 1.1005
R2748 X2.n1145 X2.n131 1.1005
R2749 X2.n1143 X2.n1142 1.1005
R2750 X2.n1141 X2.n1140 1.1005
R2751 X2.n1122 X2.n1121 1.1005
R2752 X2.n1114 X2.n152 1.1005
R2753 X2.n1127 X2.n1126 1.1005
R2754 X2.n1113 X2.n1112 1.1005
R2755 X2.n1110 X2.n152 1.1005
R2756 X2.n1108 X2.n1107 1.1005
R2757 X2.n1105 X2.n1104 1.1005
R2758 X2.n1103 X2.n156 1.1005
R2759 X2.n1100 X2.n157 1.1005
R2760 X2.n1071 X2.n1070 1.1005
R2761 X2.n1075 X2.n1068 1.1005
R2762 X2.n1077 X2.n1076 1.1005
R2763 X2.n1078 X2.n1064 1.1005
R2764 X2.n1083 X2.n1062 1.1005
R2765 X2.n1058 X2.n167 1.1005
R2766 X2.n1057 X2.n1056 1.1005
R2767 X2.n1055 X2.n168 1.1005
R2768 X2.n1046 X2.n174 1.1005
R2769 X2.n1048 X2.n1047 1.1005
R2770 X2.n1045 X2.n173 1.1005
R2771 X2.n1037 X2.n179 1.1005
R2772 X2.n1028 X2.n183 1.1005
R2773 X2.n1027 X2.n1026 1.1005
R2774 X2.n185 X2.n184 1.1005
R2775 X2.n1019 X2.n1018 1.1005
R2776 X2.n1017 X2.n188 1.1005
R2777 X2.n1016 X2.n1015 1.1005
R2778 X2.n1013 X2.n1012 1.1005
R2779 X2.n191 X2.n190 1.1005
R2780 X2.n992 X2.n991 1.1005
R2781 X2.n995 X2.n994 1.1005
R2782 X2.n987 X2.n986 1.1005
R2783 X2.n985 X2.n202 1.1005
R2784 X2.n984 X2.n983 1.1005
R2785 X2.n205 X2.n204 1.1005
R2786 X2.n969 X2.n968 1.1005
R2787 X2.n967 X2.n209 1.1005
R2788 X2.n964 X2.n210 1.1005
R2789 X2.n947 X2.n946 1.1005
R2790 X2.n951 X2.n219 1.1005
R2791 X2.n953 X2.n952 1.1005
R2792 X2.n944 X2.n218 1.1005
R2793 X2.n939 X2.n938 1.1005
R2794 X2.n927 X2.n226 1.1005
R2795 X2.n929 X2.n928 1.1005
R2796 X2.n924 X2.n923 1.1005
R2797 X2.n921 X2.n920 1.1005
R2798 X2.n917 X2.n229 1.1005
R2799 X2.n916 X2.n915 1.1005
R2800 X2.n914 X2.n230 1.1005
R2801 X2.n893 X2.n892 1.1005
R2802 X2.n889 X2.n888 1.1005
R2803 X2.n887 X2.n246 1.1005
R2804 X2.n886 X2.n885 1.1005
R2805 X2.n249 X2.n248 1.1005
R2806 X2.n878 X2.n877 1.1005
R2807 X2.n876 X2.n251 1.1005
R2808 X2.n253 X2.n252 1.1005
R2809 X2.n870 X2.n869 1.1005
R2810 X2.n867 X2.n866 1.1005
R2811 X2.n862 X2.n861 1.1005
R2812 X2.n859 X2.n858 1.1005
R2813 X2.n857 X2.n260 1.1005
R2814 X2.n851 X2.n261 1.1005
R2815 X2.n849 X2.n848 1.1005
R2816 X2.n847 X2.n264 1.1005
R2817 X2.n841 X2.n265 1.1005
R2818 X2.n840 X2.n267 1.1005
R2819 X2.n839 X2.n838 1.1005
R2820 X2.n835 X2.n834 1.1005
R2821 X2.n832 X2.n831 1.1005
R2822 X2.n825 X2.n276 1.1005
R2823 X2.n827 X2.n826 1.1005
R2824 X2.n824 X2.n275 1.1005
R2825 X2.n819 X2.n818 1.1005
R2826 X2.n382 X2.n380 1.1005
R2827 X2.n384 X2.n383 1.1005
R2828 X2.n385 X2.n374 1.1005
R2829 X2.n817 X2.n278 1.1005
R2830 X2.n816 X2.n815 1.1005
R2831 X2.n814 X2.n279 1.1005
R2832 X2.n379 X2.n280 1.1005
R2833 X2.n820 X2.n277 1.1005
R2834 X2.n823 X2.n822 1.1005
R2835 X2.n273 X2.n272 1.1005
R2836 X2.n833 X2.n271 1.1005
R2837 X2.n269 X2.n268 1.1005
R2838 X2.n843 X2.n842 1.1005
R2839 X2.n850 X2.n263 1.1005
R2840 X2.n853 X2.n852 1.1005
R2841 X2.n860 X2.n259 1.1005
R2842 X2.n257 X2.n256 1.1005
R2843 X2.n868 X2.n255 1.1005
R2844 X2.n875 X2.n874 1.1005
R2845 X2.n883 X2.n882 1.1005
R2846 X2.n884 X2.n247 1.1005
R2847 X2.n890 X2.n244 1.1005
R2848 X2.n894 X2.n891 1.1005
R2849 X2.n896 X2.n895 1.1005
R2850 X2.n897 X2.n245 1.1005
R2851 X2.n899 X2.n898 1.1005
R2852 X2.n233 X2.n232 1.1005
R2853 X2.n913 X2.n912 1.1005
R2854 X2.n919 X2.n918 1.1005
R2855 X2.n922 X2.n227 1.1005
R2856 X2.n925 X2.n225 1.1005
R2857 X2.n937 X2.n221 1.1005
R2858 X2.n936 X2.n935 1.1005
R2859 X2.n934 X2.n222 1.1005
R2860 X2.n926 X2.n223 1.1005
R2861 X2.n940 X2.n220 1.1005
R2862 X2.n943 X2.n942 1.1005
R2863 X2.n950 X2.n949 1.1005
R2864 X2.n945 X2.n211 1.1005
R2865 X2.n966 X2.n965 1.1005
R2866 X2.n975 X2.n974 1.1005
R2867 X2.n973 X2.n207 1.1005
R2868 X2.n972 X2.n971 1.1005
R2869 X2.n970 X2.n208 1.1005
R2870 X2.n981 X2.n980 1.1005
R2871 X2.n982 X2.n203 1.1005
R2872 X2.n988 X2.n200 1.1005
R2873 X2.n993 X2.n201 1.1005
R2874 X2.n990 X2.n989 1.1005
R2875 X2.n1014 X2.n189 1.1005
R2876 X2.n1020 X2.n187 1.1005
R2877 X2.n1022 X2.n1021 1.1005
R2878 X2.n1030 X2.n1029 1.1005
R2879 X2.n1039 X2.n1038 1.1005
R2880 X2.n1036 X2.n178 1.1005
R2881 X2.n1035 X2.n1034 1.1005
R2882 X2.n181 X2.n180 1.1005
R2883 X2.n176 X2.n175 1.1005
R2884 X2.n1044 X2.n1043 1.1005
R2885 X2.n171 X2.n170 1.1005
R2886 X2.n1054 X2.n1053 1.1005
R2887 X2.n1060 X2.n1059 1.1005
R2888 X2.n1085 X2.n1084 1.1005
R2889 X2.n1086 X2.n166 1.1005
R2890 X2.n1088 X2.n1087 1.1005
R2891 X2.n1061 X2.n165 1.1005
R2892 X2.n1082 X2.n1081 1.1005
R2893 X2.n1080 X2.n1079 1.1005
R2894 X2.n1074 X2.n1073 1.1005
R2895 X2.n1069 X2.n158 1.1005
R2896 X2.n1102 X2.n1101 1.1005
R2897 X2.n1112 X2.n1111 1.1005
R2898 X2.n1106 X2.n155 1.1005
R2899 X2.n1109 X2.n151 1.1005
R2900 X2.n390 X2.n372 1.1005
R2901 X2.n401 X2.n400 1.1005
R2902 X2.n423 X2.n365 1.1005
R2903 X2.n470 X2.n469 1.1005
R2904 X2.n490 X2.n489 1.1005
R2905 X2.n511 X2.n334 1.1005
R2906 X2.n378 X2.n375 1.1005
R2907 X2.n387 X2.n373 1.1005
R2908 X2.n392 X2.n391 1.1005
R2909 X2.n731 X2.n730 1.1005
R2910 X2.n737 X2.n736 1.1005
R2911 X2.n532 X2.n531 1.1005
R2912 X2.n750 X2.n749 1.1005
R2913 X2.n516 X2.n319 1.1005
R2914 X2.n513 X2.n512 1.1005
R2915 X2.n499 X2.n498 1.1005
R2916 X2.n488 X2.n339 1.1005
R2917 X2.n479 X2.n478 1.1005
R2918 X2.n468 X2.n348 1.1005
R2919 X2.n461 X2.n460 1.1005
R2920 X2.n441 X2.n440 1.1005
R2921 X2.n425 X2.n424 1.1005
R2922 X2.n413 X2.n412 1.1005
R2923 X2.n399 X2.n370 1.1005
R2924 X2.n389 X2.n388 1.1005
R2925 X2.n376 X2.n375 1.1005
R2926 X2.n387 X2.n386 1.1005
R2927 X2.n1320 X2.n1319 0.733833
R2928 X2.n1128 X2.n1127 0.733833
R2929 X2.n388 X2.n285 0.733833
R2930 X2.n727 X2.n726 0.733833
R2931 X2.n502 X2.n334 0.573769
R2932 X2.n419 X2.n365 0.573769
R2933 X2.n491 X2.n490 0.573695
R2934 X2.n402 X2.n401 0.573695
R2935 X2.n469 X2.n349 0.573346
R2936 X2.n480 X2.n346 0.573297
R2937 X2.n154 X2.n152 0.550549
R2938 X2.n387 X2.n377 0.550549
R2939 X2.n513 X2.n333 0.39244
R2940 X2.n425 X2.n364 0.39244
R2941 X2.n486 X2.n339 0.389994
R2942 X2.n395 X2.n370 0.389994
R2943 X2.n351 X2.n348 0.387191
R2944 X2.n751 X2.n521 0.384705
R2945 X2.n448 X2.n354 0.384705
R2946 X2.n514 X2.n332 0.384705
R2947 X2.n427 X2.n426 0.384705
R2948 X2.n752 X2.n321 0.382331
R2949 X2.n442 X2.n357 0.382331
R2950 X2.n515 X2.n322 0.382034
R2951 X2.n360 X2.n359 0.382034
R2952 X2.n500 X2.n335 0.379547
R2953 X2.n463 X2.n462 0.379547
R2954 X2.n414 X2.n366 0.379547
R2955 X2.n500 X2.n338 0.375976
R2956 X2.n414 X2.n369 0.375976
R2957 X2.n462 X2.n353 0.375884
R2958 X2.n515 X2.n326 0.374982
R2959 X2.n432 X2.n359 0.374982
R2960 X2.n753 X2.n752 0.374889
R2961 X2.n443 X2.n442 0.374889
R2962 X2.n751 X2.n522 0.373984
R2963 X2.n355 X2.n354 0.373984
R2964 X2.n514 X2.n327 0.373891
R2965 X2.n426 X2.n363 0.373891
R2966 X2.n481 X2.n480 0.280767
R2967 X2.n728 X2.n727 0.275034
R2968 X2.n3 X2.n2 0.182739
R2969 X2 X2.n1377 0.103107
R2970 X2 X2.n1378 0.08058
R2971 X2.n2 X2 0.0563209
R2972 X2.n4 X2 0.0445
R2973 X2.n1363 X2.n1362 0.0405
R2974 X2.n1362 X2.n1361 0.0405
R2975 X2.n1361 X2.n21 0.0405
R2976 X2.n1357 X2.n21 0.0405
R2977 X2.n1357 X2.n1356 0.0405
R2978 X2.n1356 X2.n1355 0.0405
R2979 X2.n1355 X2.n26 0.0405
R2980 X2.n1351 X2.n26 0.0405
R2981 X2.n1351 X2.n1350 0.0405
R2982 X2.n1350 X2.n1349 0.0405
R2983 X2.n1349 X2.n31 0.0405
R2984 X2.n1345 X2.n31 0.0405
R2985 X2.n1345 X2.n1344 0.0405
R2986 X2.n1344 X2.n1343 0.0405
R2987 X2.n1339 X2.n36 0.0405
R2988 X2.n1339 X2.n1338 0.0405
R2989 X2.n1338 X2.n1337 0.0405
R2990 X2.n1337 X2.n41 0.0405
R2991 X2.n1333 X2.n41 0.0405
R2992 X2.n1333 X2.n1332 0.0405
R2993 X2.n1332 X2.n1331 0.0405
R2994 X2.n1331 X2.n46 0.0405
R2995 X2.n1327 X2.n46 0.0405
R2996 X2.n1327 X2.n1326 0.0405
R2997 X2.n1326 X2.n1325 0.0405
R2998 X2.n1325 X2.n51 0.0405
R2999 X2.n1364 X2.n17 0.0405
R3000 X2.n1360 X2.n17 0.0405
R3001 X2.n1360 X2.n1359 0.0405
R3002 X2.n1359 X2.n1358 0.0405
R3003 X2.n1358 X2.n22 0.0405
R3004 X2.n1354 X2.n22 0.0405
R3005 X2.n1354 X2.n1353 0.0405
R3006 X2.n1353 X2.n1352 0.0405
R3007 X2.n1352 X2.n27 0.0405
R3008 X2.n1348 X2.n27 0.0405
R3009 X2.n1348 X2.n1347 0.0405
R3010 X2.n1347 X2.n1346 0.0405
R3011 X2.n1346 X2.n32 0.0405
R3012 X2.n1342 X2.n32 0.0405
R3013 X2.n1341 X2.n1340 0.0405
R3014 X2.n1340 X2.n37 0.0405
R3015 X2.n1336 X2.n37 0.0405
R3016 X2.n1336 X2.n1335 0.0405
R3017 X2.n1335 X2.n1334 0.0405
R3018 X2.n1334 X2.n42 0.0405
R3019 X2.n1330 X2.n42 0.0405
R3020 X2.n1330 X2.n1329 0.0405
R3021 X2.n1329 X2.n1328 0.0405
R3022 X2.n1328 X2.n47 0.0405
R3023 X2.n1324 X2.n47 0.0405
R3024 X2.n1324 X2.n1323 0.0405
R3025 X2.n810 X2.n282 0.0405
R3026 X2.n810 X2.n283 0.0405
R3027 X2.n806 X2.n283 0.0405
R3028 X2.n806 X2.n805 0.0405
R3029 X2.n805 X2.n804 0.0405
R3030 X2.n804 X2.n801 0.0405
R3031 X2.n801 X2.n240 0.0405
R3032 X2.n903 X2.n240 0.0405
R3033 X2.n903 X2.n235 0.0405
R3034 X2.n908 X2.n235 0.0405
R3035 X2.n908 X2.n238 0.0405
R3036 X2.n238 X2.n215 0.0405
R3037 X2.n956 X2.n215 0.0405
R3038 X2.n956 X2.n213 0.0405
R3039 X2.n960 X2.n196 0.0405
R3040 X2.n999 X2.n196 0.0405
R3041 X2.n999 X2.n193 0.0405
R3042 X2.n1008 X2.n193 0.0405
R3043 X2.n1008 X2.n194 0.0405
R3044 X2.n1004 X2.n194 0.0405
R3045 X2.n1004 X2.n1003 0.0405
R3046 X2.n1003 X2.n162 0.0405
R3047 X2.n1091 X2.n162 0.0405
R3048 X2.n1091 X2.n160 0.0405
R3049 X2.n1095 X2.n160 0.0405
R3050 X2.n1095 X2.n148 0.0405
R3051 X2.n809 X2.n799 0.0405
R3052 X2.n809 X2.n808 0.0405
R3053 X2.n808 X2.n807 0.0405
R3054 X2.n807 X2.n800 0.0405
R3055 X2.n803 X2.n800 0.0405
R3056 X2.n803 X2.n802 0.0405
R3057 X2.n802 X2.n239 0.0405
R3058 X2.n904 X2.n239 0.0405
R3059 X2.n905 X2.n904 0.0405
R3060 X2.n907 X2.n905 0.0405
R3061 X2.n907 X2.n906 0.0405
R3062 X2.n906 X2.n214 0.0405
R3063 X2.n957 X2.n214 0.0405
R3064 X2.n958 X2.n957 0.0405
R3065 X2.n959 X2.n195 0.0405
R3066 X2.n1000 X2.n195 0.0405
R3067 X2.n1001 X2.n1000 0.0405
R3068 X2.n1007 X2.n1001 0.0405
R3069 X2.n1007 X2.n1006 0.0405
R3070 X2.n1006 X2.n1005 0.0405
R3071 X2.n1005 X2.n1002 0.0405
R3072 X2.n1002 X2.n161 0.0405
R3073 X2.n1092 X2.n161 0.0405
R3074 X2.n1093 X2.n1092 0.0405
R3075 X2.n1094 X2.n1093 0.0405
R3076 X2.n1094 X2.n147 0.0405
R3077 X2.n1343 X2.n36 0.0360676
R3078 X2.n1342 X2.n1341 0.0360676
R3079 X2.n960 X2.n213 0.0360676
R3080 X2.n959 X2.n958 0.0360676
R3081 X2.n1132 X2.n1131 0.0360676
R3082 X2.n1132 X2.n137 0.0360676
R3083 X2.n1152 X2.n137 0.0360676
R3084 X2.n1153 X2.n1152 0.0360676
R3085 X2.n1154 X2.n1153 0.0360676
R3086 X2.n1154 X2.n123 0.0360676
R3087 X2.n1175 X2.n123 0.0360676
R3088 X2.n1176 X2.n1175 0.0360676
R3089 X2.n1177 X2.n1176 0.0360676
R3090 X2.n1178 X2.n1177 0.0360676
R3091 X2.n1178 X2.n111 0.0360676
R3092 X2.n1206 X2.n111 0.0360676
R3093 X2.n1207 X2.n1206 0.0360676
R3094 X2.n1208 X2.n1207 0.0360676
R3095 X2.n1209 X2.n1208 0.0360676
R3096 X2.n1209 X2.n94 0.0360676
R3097 X2.n1230 X2.n94 0.0360676
R3098 X2.n1231 X2.n1230 0.0360676
R3099 X2.n1232 X2.n1231 0.0360676
R3100 X2.n1232 X2.n84 0.0360676
R3101 X2.n1253 X2.n84 0.0360676
R3102 X2.n1254 X2.n1253 0.0360676
R3103 X2.n1255 X2.n1254 0.0360676
R3104 X2.n1256 X2.n1255 0.0360676
R3105 X2.n1256 X2.n73 0.0360676
R3106 X2.n1284 X2.n73 0.0360676
R3107 X2.n1285 X2.n1284 0.0360676
R3108 X2.n1286 X2.n1285 0.0360676
R3109 X2.n1286 X2.n64 0.0360676
R3110 X2.n1308 X2.n64 0.0360676
R3111 X2.n1309 X2.n1308 0.0360676
R3112 X2.n1310 X2.n1309 0.0360676
R3113 X2.n1310 X2.n52 0.0360676
R3114 X2.n1133 X2.n146 0.0360676
R3115 X2.n1133 X2.n138 0.0360676
R3116 X2.n1151 X2.n138 0.0360676
R3117 X2.n1151 X2.n136 0.0360676
R3118 X2.n1155 X2.n136 0.0360676
R3119 X2.n1155 X2.n124 0.0360676
R3120 X2.n1174 X2.n124 0.0360676
R3121 X2.n1174 X2.n122 0.0360676
R3122 X2.n1180 X2.n122 0.0360676
R3123 X2.n1180 X2.n1179 0.0360676
R3124 X2.n1179 X2.n112 0.0360676
R3125 X2.n1205 X2.n112 0.0360676
R3126 X2.n1205 X2.n110 0.0360676
R3127 X2.n1211 X2.n110 0.0360676
R3128 X2.n1211 X2.n1210 0.0360676
R3129 X2.n1210 X2.n95 0.0360676
R3130 X2.n1229 X2.n95 0.0360676
R3131 X2.n1229 X2.n93 0.0360676
R3132 X2.n1233 X2.n93 0.0360676
R3133 X2.n1233 X2.n85 0.0360676
R3134 X2.n1252 X2.n85 0.0360676
R3135 X2.n1252 X2.n83 0.0360676
R3136 X2.n1258 X2.n83 0.0360676
R3137 X2.n1258 X2.n1257 0.0360676
R3138 X2.n1257 X2.n74 0.0360676
R3139 X2.n1283 X2.n74 0.0360676
R3140 X2.n1283 X2.n72 0.0360676
R3141 X2.n1287 X2.n72 0.0360676
R3142 X2.n1287 X2.n65 0.0360676
R3143 X2.n1307 X2.n65 0.0360676
R3144 X2.n1307 X2.n63 0.0360676
R3145 X2.n1311 X2.n63 0.0360676
R3146 X2.n1311 X2.n53 0.0360676
R3147 X2.n796 X2.n795 0.0360676
R3148 X2.n795 X2.n288 0.0360676
R3149 X2.n791 X2.n288 0.0360676
R3150 X2.n791 X2.n790 0.0360676
R3151 X2.n790 X2.n789 0.0360676
R3152 X2.n789 X2.n293 0.0360676
R3153 X2.n785 X2.n293 0.0360676
R3154 X2.n785 X2.n784 0.0360676
R3155 X2.n784 X2.n783 0.0360676
R3156 X2.n783 X2.n298 0.0360676
R3157 X2.n779 X2.n298 0.0360676
R3158 X2.n779 X2.n778 0.0360676
R3159 X2.n778 X2.n777 0.0360676
R3160 X2.n777 X2.n303 0.0360676
R3161 X2.n773 X2.n303 0.0360676
R3162 X2.n773 X2.n772 0.0360676
R3163 X2.n772 X2.n771 0.0360676
R3164 X2.n771 X2.n308 0.0360676
R3165 X2.n767 X2.n308 0.0360676
R3166 X2.n767 X2.n766 0.0360676
R3167 X2.n766 X2.n765 0.0360676
R3168 X2.n765 X2.n313 0.0360676
R3169 X2.n761 X2.n313 0.0360676
R3170 X2.n761 X2.n760 0.0360676
R3171 X2.n760 X2.n759 0.0360676
R3172 X2.n759 X2.n7 0.0360676
R3173 X2.n1375 X2.n7 0.0360676
R3174 X2.n1375 X2.n1374 0.0360676
R3175 X2.n1374 X2.n1373 0.0360676
R3176 X2.n1373 X2.n11 0.0360676
R3177 X2.n1369 X2.n11 0.0360676
R3178 X2.n1369 X2.n1368 0.0360676
R3179 X2.n1368 X2.n1367 0.0360676
R3180 X2.n794 X2.n284 0.0360676
R3181 X2.n794 X2.n793 0.0360676
R3182 X2.n793 X2.n792 0.0360676
R3183 X2.n792 X2.n289 0.0360676
R3184 X2.n788 X2.n289 0.0360676
R3185 X2.n788 X2.n787 0.0360676
R3186 X2.n787 X2.n786 0.0360676
R3187 X2.n786 X2.n294 0.0360676
R3188 X2.n782 X2.n294 0.0360676
R3189 X2.n782 X2.n781 0.0360676
R3190 X2.n781 X2.n780 0.0360676
R3191 X2.n780 X2.n299 0.0360676
R3192 X2.n776 X2.n299 0.0360676
R3193 X2.n776 X2.n775 0.0360676
R3194 X2.n775 X2.n774 0.0360676
R3195 X2.n774 X2.n304 0.0360676
R3196 X2.n770 X2.n304 0.0360676
R3197 X2.n770 X2.n769 0.0360676
R3198 X2.n769 X2.n768 0.0360676
R3199 X2.n768 X2.n309 0.0360676
R3200 X2.n764 X2.n309 0.0360676
R3201 X2.n764 X2.n763 0.0360676
R3202 X2.n763 X2.n762 0.0360676
R3203 X2.n762 X2.n314 0.0360676
R3204 X2.n758 X2.n314 0.0360676
R3205 X2.n758 X2.n5 0.0360676
R3206 X2.n1376 X2.n6 0.0360676
R3207 X2.n1372 X2.n6 0.0360676
R3208 X2.n1372 X2.n1371 0.0360676
R3209 X2.n1371 X2.n1370 0.0360676
R3210 X2.n1370 X2.n12 0.0360676
R3211 X2.n1366 X2.n12 0.0360676
R3212 X2.n1363 X2.n16 0.0234189
R3213 X2.n1365 X2.n1364 0.0234189
R3214 X2.n797 X2.n282 0.0234189
R3215 X2.n799 X2.n798 0.0234189
R3216 X2.n1321 X2.n51 0.0233108
R3217 X2.n1323 X2.n1322 0.0233108
R3218 X2.n1129 X2.n148 0.0233108
R3219 X2.n1130 X2.n147 0.0233108
R3220 X2.n1377 X2.n5 0.0228784
R3221 X2.n1131 X2.n1130 0.0227703
R3222 X2.n1129 X2.n146 0.0227703
R3223 X2.n797 X2.n796 0.0227703
R3224 X2.n798 X2.n284 0.0227703
R3225 X2.n717 X2.n716 0.0188784
R3226 X2.n713 X2.n712 0.0188784
R3227 X2.n709 X2.n708 0.0188784
R3228 X2.n705 X2.n704 0.0188784
R3229 X2.n560 X2.n559 0.0188784
R3230 X2.n690 X2.n563 0.0188784
R3231 X2.n568 X2.n567 0.0188784
R3232 X2.n684 X2.n683 0.0188784
R3233 X2.n679 X2.n678 0.0188784
R3234 X2.n676 X2.n571 0.0188784
R3235 X2.n669 X2.n667 0.0188784
R3236 X2.n664 X2.n663 0.0188784
R3237 X2.n660 X2.n659 0.0188784
R3238 X2.n656 X2.n655 0.0188784
R3239 X2.n652 X2.n651 0.0188784
R3240 X2.n583 X2.n582 0.0188784
R3241 X2.n644 X2.n643 0.0188784
R3242 X2.n641 X2.n586 0.0188784
R3243 X2.n631 X2.n630 0.0188784
R3244 X2.n626 X2.n625 0.0188784
R3245 X2.n623 X2.n594 0.0188784
R3246 X2.n616 X2.n615 0.0188784
R3247 X2.n613 X2.n612 0.0188784
R3248 X2.n829 X2.n828 0.0188784
R3249 X2.n837 X2.n836 0.0188784
R3250 X2.n846 X2.n845 0.0188784
R3251 X2.n856 X2.n855 0.0188784
R3252 X2.n865 X2.n864 0.0188784
R3253 X2.n880 X2.n241 0.0188784
R3254 X2.n901 X2.n243 0.0188784
R3255 X2.n910 X2.n234 0.0188784
R3256 X2.n236 X2.n231 0.0188784
R3257 X2.n930 X2.n224 0.0188784
R3258 X2.n933 X2.n932 0.0188784
R3259 X2.n954 X2.n217 0.0188784
R3260 X2.n963 X2.n962 0.0188784
R3261 X2.n976 X2.n206 0.0188784
R3262 X2.n978 X2.n197 0.0188784
R3263 X2.n997 X2.n199 0.0188784
R3264 X2.n1010 X2.n192 0.0188784
R3265 X2.n1024 X2.n186 0.0188784
R3266 X2.n1041 X2.n1040 0.0188784
R3267 X2.n1051 X2.n1049 0.0188784
R3268 X2.n169 X2.n163 0.0188784
R3269 X2.n1089 X2.n164 0.0188784
R3270 X2.n1067 X2.n1066 0.0188784
R3271 X2.n1128 X2.n150 0.0188784
R3272 X2.n1118 X2.n145 0.0188784
R3273 X2.n1138 X2.n1135 0.0188784
R3274 X2.n1136 X2.n139 0.0188784
R3275 X2.n1221 X2.n96 0.0188784
R3276 X2.n1227 X2.n97 0.0188784
R3277 X2.n102 X2.n92 0.0188784
R3278 X2.n1237 X2.n1235 0.0188784
R3279 X2.n393 X2.n285 0.0188784
R3280 X2.n397 X2.n396 0.0188784
R3281 X2.n410 X2.n405 0.0188784
R3282 X2.n408 X2.n407 0.0188784
R3283 X2.n484 X2.n483 0.0188784
R3284 X2.n493 X2.n345 0.0188784
R3285 X2.n496 X2.n495 0.0188784
R3286 X2.n343 X2.n342 0.0188784
R3287 X2.n722 X2.n721 0.0187703
R3288 X2.n718 X2.n717 0.0187703
R3289 X2.n697 X2.n696 0.0187703
R3290 X2.n694 X2.n563 0.0187703
R3291 X2.n669 X2.n668 0.0187703
R3292 X2.n637 X2.n586 0.0187703
R3293 X2.n591 X2.n590 0.0187703
R3294 X2.n612 X2.n599 0.0187703
R3295 X2.n608 X2.n607 0.0187703
R3296 X2.n813 X2.n812 0.0187703
R3297 X2.n828 X2.n274 0.0187703
R3298 X2.n872 X2.n871 0.0187703
R3299 X2.n880 X2.n879 0.0187703
R3300 X2.n932 X2.n216 0.0187703
R3301 X2.n1025 X2.n1024 0.0187703
R3302 X2.n1033 X2.n1032 0.0187703
R3303 X2.n1067 X2.n159 0.0187703
R3304 X2.n1099 X2.n1098 0.0187703
R3305 X2.n1146 X2.n135 0.0187703
R3306 X2.n1160 X2.n1157 0.0187703
R3307 X2.n1158 X2.n125 0.0187703
R3308 X2.n1172 X2.n126 0.0187703
R3309 X2.n129 X2.n121 0.0187703
R3310 X2.n1183 X2.n1182 0.0187703
R3311 X2.n1188 X2.n1187 0.0187703
R3312 X2.n1190 X2.n113 0.0187703
R3313 X2.n1203 X2.n114 0.0187703
R3314 X2.n1195 X2.n109 0.0187703
R3315 X2.n1214 X2.n1213 0.0187703
R3316 X2.n1219 X2.n1218 0.0187703
R3317 X2.n1250 X2.n87 0.0187703
R3318 X2.n1242 X2.n82 0.0187703
R3319 X2.n1261 X2.n1260 0.0187703
R3320 X2.n1266 X2.n1265 0.0187703
R3321 X2.n1268 X2.n75 0.0187703
R3322 X2.n1281 X2.n76 0.0187703
R3323 X2.n1277 X2.n71 0.0187703
R3324 X2.n1292 X2.n1289 0.0187703
R3325 X2.n1290 X2.n66 0.0187703
R3326 X2.n1305 X2.n67 0.0187703
R3327 X2.n1300 X2.n62 0.0187703
R3328 X2.n1314 X2.n1313 0.0187703
R3329 X2.n421 X2.n420 0.0187703
R3330 X2.n417 X2.n416 0.0187703
R3331 X2.n430 X2.n429 0.0187703
R3332 X2.n435 X2.n434 0.0187703
R3333 X2.n438 X2.n437 0.0187703
R3334 X2.n446 X2.n445 0.0187703
R3335 X2.n451 X2.n450 0.0187703
R3336 X2.n458 X2.n457 0.0187703
R3337 X2.n455 X2.n454 0.0187703
R3338 X2.n466 X2.n465 0.0187703
R3339 X2.n473 X2.n472 0.0187703
R3340 X2.n476 X2.n475 0.0187703
R3341 X2.n509 X2.n503 0.0187703
R3342 X2.n507 X2.n505 0.0187703
R3343 X2.n330 X2.n329 0.0187703
R3344 X2.n324 X2.n317 0.0187703
R3345 X2.n756 X2.n318 0.0187703
R3346 X2.n519 X2.n518 0.0187703
R3347 X2.n526 X2.n525 0.0187703
R3348 X2.n747 X2.n746 0.0187703
R3349 X2.n744 X2.n743 0.0187703
R3350 X2.n537 X2.n536 0.0187703
R3351 X2.n734 X2.n733 0.0187703
R3352 X2.n542 X2.n541 0.0187703
R3353 X2.n713 X2.n20 0.0185541
R3354 X2.n616 X2.n49 0.0185541
R3355 X2.n836 X2.n270 0.0185541
R3356 X2.n1065 X2.n164 0.0185541
R3357 X2.n1149 X2.n140 0.0184459
R3358 X2.n1251 X2.n86 0.0184459
R3359 X2.n367 X2.n291 0.0184459
R3360 X2.n336 X2.n312 0.0184459
R3361 X2.n664 X2.n34 0.0182297
R3362 X2.n955 X2.n954 0.0182297
R3363 X2.n1150 X2.n1149 0.0181216
R3364 X2.n1236 X2.n86 0.0181216
R3365 X2.n367 X2.n290 0.0181216
R3366 X2.n336 X2.n311 0.0181216
R3367 X2.n696 X2.n695 0.0175811
R3368 X2.n590 X2.n43 0.0175811
R3369 X2.n872 X2.n250 0.0175811
R3370 X2.n1032 X2.n182 0.0175811
R3371 X2.n1156 X2.n135 0.0173649
R3372 X2.n1241 X2.n87 0.0173649
R3373 X2.n421 X2.n292 0.0173649
R3374 X2.n509 X2.n508 0.0173649
R3375 X2.n1137 X2.n1136 0.0170405
R3376 X2.n1235 X2.n1234 0.0170405
R3377 X2.n409 X2.n408 0.0170405
R3378 X2.n343 X2.n310 0.0170405
R3379 X2.n567 X2.n28 0.0167162
R3380 X2.n643 X2.n642 0.0167162
R3381 X2.n902 X2.n901 0.0167162
R3382 X2.n1010 X2.n1009 0.0167162
R3383 X2.n1160 X2.n1159 0.0162838
R3384 X2.n1259 X2.n82 0.0162838
R3385 X2.n416 X2.n361 0.0162838
R3386 X2.n505 X2.n315 0.0162838
R3387 X2.n571 X2.n33 0.0159595
R3388 X2.n656 X2.n576 0.0159595
R3389 X2.n931 X2.n930 0.0159595
R3390 X2.n961 X2.n206 0.0159595
R3391 X2.n1135 X2.n1134 0.0159595
R3392 X2.n102 X2.n101 0.0159595
R3393 X2.n405 X2.n287 0.0159595
R3394 X2.n495 X2.n494 0.0159595
R3395 X2.n721 X2.n19 0.0157432
R3396 X2.n608 X2.n50 0.0157432
R3397 X2.n812 X2.n811 0.0157432
R3398 X2.n1099 X2.n1096 0.0157432
R3399 X2.n709 X2.n551 0.0152027
R3400 X2.n594 X2.n48 0.0152027
R3401 X2.n845 X2.n266 0.0152027
R3402 X2.n1090 X2.n163 0.0152027
R3403 X2.n1173 X2.n125 0.0152027
R3404 X2.n1261 X2.n80 0.0152027
R3405 X2.n430 X2.n295 0.0152027
R3406 X2.n329 X2.n316 0.0152027
R3407 X2.n660 X2.n35 0.0148784
R3408 X2.n963 X2.n212 0.0148784
R3409 X2.n1118 X2.n1117 0.0148784
R3410 X2.n1228 X2.n1227 0.0148784
R3411 X2.n397 X2.n286 0.0148784
R3412 X2.n345 X2.n307 0.0148784
R3413 X2.n560 X2.n25 0.0141216
R3414 X2.n631 X2.n44 0.0141216
R3415 X2.n865 X2.n254 0.0141216
R3416 X2.n1040 X2.n177 0.0141216
R3417 X2.n128 X2.n126 0.0141216
R3418 X2.n1267 X2.n1266 0.0141216
R3419 X2.n435 X2.n296 0.0141216
R3420 X2.n757 X2.n317 0.0141216
R3421 X2.n1322 X2.n52 0.0137973
R3422 X2.n1321 X2.n53 0.0137973
R3423 X2.n1221 X2.n1220 0.0137973
R3424 X2.n1320 X2.n55 0.0137973
R3425 X2.n483 X2.n306 0.0137973
R3426 X2.n726 X2.n15 0.0137973
R3427 X2.n1367 X2.n16 0.0137973
R3428 X2.n1366 X2.n1365 0.0137973
R3429 X2.n1377 X2.n1376 0.0136892
R3430 X2.n1318 X2.n1317 0.0134381
R3431 X2.n684 X2.n29 0.0133649
R3432 X2.n583 X2.n40 0.0133649
R3433 X2.n242 X2.n234 0.0133649
R3434 X2.n199 X2.n198 0.0133649
R3435 X2.n1181 X2.n121 0.0130405
R3436 X2.n1282 X2.n75 0.0130405
R3437 X2.n437 X2.n297 0.0130405
R3438 X2.n517 X2.n318 0.0130405
R3439 X2.n1218 X2.n107 0.0128243
R3440 X2.n1314 X2.n1312 0.0128243
R3441 X2.n476 X2.n305 0.0128243
R3442 X2.n541 X2.n14 0.0128243
R3443 X2.n678 X2.n677 0.0126081
R3444 X2.n652 X2.n38 0.0126081
R3445 X2.n237 X2.n236 0.0126081
R3446 X2.n978 X2.n977 0.0126081
R3447 X2.n725 X2.n18 0.0123919
R3448 X2.n605 X2.n54 0.0123919
R3449 X2.n381 X2.n281 0.0123919
R3450 X2.n1097 X2.n149 0.0123919
R3451 X2.n1183 X2.n119 0.0119595
R3452 X2.n1276 X2.n76 0.0119595
R3453 X2.n446 X2.n356 0.0119595
R3454 X2.n519 X2.n8 0.0119595
R3455 X2.n705 X2.n23 0.0118514
R3456 X2.n625 X2.n624 0.0118514
R3457 X2.n855 X2.n262 0.0118514
R3458 X2.n1051 X2.n1050 0.0118514
R3459 X2.n1213 X2.n1212 0.0117432
R3460 X2.n1300 X2.n1299 0.0117432
R3461 X2.n472 X2.n350 0.0117432
R3462 X2.n734 X2.n13 0.0117432
R3463 X2.n728 X2.n545 0.0116588
R3464 X2.n726 X2.n725 0.011527
R3465 X2.n381 X2.n285 0.011527
R3466 X2.n1320 X2.n54 0.0114189
R3467 X2.n1128 X2.n149 0.0114189
R3468 X2.n414 X2.n413 0.0109762
R3469 X2.n426 X2.n425 0.0109762
R3470 X2.n441 X2.n359 0.0109762
R3471 X2.n442 X2.n354 0.0109762
R3472 X2.n462 X2.n461 0.0109762
R3473 X2.n479 X2.n348 0.0109762
R3474 X2.n480 X2.n339 0.0109762
R3475 X2.n500 X2.n499 0.0109762
R3476 X2.n514 X2.n513 0.0109762
R3477 X2.n516 X2.n515 0.0109762
R3478 X2.n752 X2.n751 0.0109762
R3479 X2.n555 X2.n554 0.0109762
R3480 X2.n556 X2.n555 0.0109762
R3481 X2.n557 X2.n556 0.0109762
R3482 X2.n701 X2.n557 0.0109762
R3483 X2.n701 X2.n700 0.0109762
R3484 X2.n700 X2.n558 0.0109762
R3485 X2.n688 X2.n558 0.0109762
R3486 X2.n688 X2.n687 0.0109762
R3487 X2.n687 X2.n566 0.0109762
R3488 X2.n673 X2.n566 0.0109762
R3489 X2.n673 X2.n672 0.0109762
R3490 X2.n579 X2.n573 0.0109762
R3491 X2.n580 X2.n579 0.0109762
R3492 X2.n648 X2.n580 0.0109762
R3493 X2.n648 X2.n647 0.0109762
R3494 X2.n647 X2.n581 0.0109762
R3495 X2.n635 X2.n581 0.0109762
R3496 X2.n635 X2.n634 0.0109762
R3497 X2.n634 X2.n589 0.0109762
R3498 X2.n620 X2.n589 0.0109762
R3499 X2.n620 X2.n619 0.0109762
R3500 X2.n619 X2.n596 0.0109762
R3501 X2.n603 X2.n596 0.0109762
R3502 X2.n1142 X2.n1141 0.0109762
R3503 X2.n1163 X2.n131 0.0109762
R3504 X2.n1168 X2.n1164 0.0109762
R3505 X2.n1167 X2.n117 0.0109762
R3506 X2.n1200 X2.n1193 0.0109762
R3507 X2.n1199 X2.n105 0.0109762
R3508 X2.n1224 X2.n1223 0.0109762
R3509 X2.n1240 X2.n90 0.0109762
R3510 X2.n1247 X2.n1246 0.0109762
R3511 X2.n1271 X2.n78 0.0109762
R3512 X2.n1272 X2.n69 0.0109762
R3513 X2.n1296 X2.n1295 0.0109762
R3514 X2.n1317 X2.n60 0.0109762
R3515 X2.n413 X2.n370 0.01095
R3516 X2.n425 X2.n414 0.01095
R3517 X2.n426 X2.n359 0.01095
R3518 X2.n442 X2.n441 0.01095
R3519 X2.n461 X2.n354 0.01095
R3520 X2.n462 X2.n348 0.01095
R3521 X2.n480 X2.n479 0.01095
R3522 X2.n499 X2.n339 0.01095
R3523 X2.n513 X2.n500 0.01095
R3524 X2.n515 X2.n514 0.01095
R3525 X2.n752 X2.n516 0.01095
R3526 X2.n751 X2.n750 0.01095
R3527 X2.n672 X2.n573 0.01095
R3528 X2.n603 X2.n602 0.01095
R3529 X2.n1142 X2.n131 0.01095
R3530 X2.n1164 X2.n1163 0.01095
R3531 X2.n1168 X2.n1167 0.01095
R3532 X2.n1193 X2.n117 0.01095
R3533 X2.n1200 X2.n1199 0.01095
R3534 X2.n1223 X2.n105 0.01095
R3535 X2.n1224 X2.n90 0.01095
R3536 X2.n1247 X2.n1240 0.01095
R3537 X2.n1246 X2.n78 0.01095
R3538 X2.n1272 X2.n1271 0.01095
R3539 X2.n1295 X2.n69 0.01095
R3540 X2.n1296 X2.n60 0.01095
R3541 X2.n1189 X2.n1188 0.0108784
R3542 X2.n1288 X2.n71 0.0108784
R3543 X2.n451 X2.n300 0.0108784
R3544 X2.n526 X2.n9 0.0108784
R3545 X2.n704 X2.n24 0.0107703
R3546 X2.n626 X2.n45 0.0107703
R3547 X2.n856 X2.n258 0.0107703
R3548 X2.n1049 X2.n172 0.0107703
R3549 X2.n1195 X2.n1194 0.0106622
R3550 X2.n1306 X2.n1305 0.0106622
R3551 X2.n465 X2.n302 0.0106622
R3552 X2.n536 X2.n530 0.0106622
R3553 X2.n554 X2.n545 0.0106095
R3554 X2.n679 X2.n30 0.0100135
R3555 X2.n651 X2.n39 0.0100135
R3556 X2.n909 X2.n231 0.0100135
R3557 X2.n998 X2.n197 0.0100135
R3558 X2.n1204 X2.n113 0.0097973
R3559 X2.n1292 X2.n1291 0.0097973
R3560 X2.n458 X2.n301 0.0097973
R3561 X2.n747 X2.n10 0.0097973
R3562 X2.n729 X2.n728 0.00967266
R3563 X2.n1204 X2.n1203 0.00958108
R3564 X2.n1291 X2.n1290 0.00958108
R3565 X2.n455 X2.n301 0.00958108
R3566 X2.n744 X2.n10 0.00958108
R3567 X2.n683 X2.n30 0.00925676
R3568 X2.n582 X2.n39 0.00925676
R3569 X2.n910 X2.n909 0.00925676
R3570 X2.n998 X2.n997 0.00925676
R3571 X2.n469 X2.n348 0.00880612
R3572 X2.n1194 X2.n114 0.00871622
R3573 X2.n1306 X2.n66 0.00871622
R3574 X2.n454 X2.n302 0.00871622
R3575 X2.n743 X2.n530 0.00871622
R3576 X2.n559 X2.n24 0.0085
R3577 X2.n630 X2.n45 0.0085
R3578 X2.n864 X2.n258 0.0085
R3579 X2.n1041 X2.n172 0.0085
R3580 X2.n1190 X2.n1189 0.0085
R3581 X2.n1289 X2.n1288 0.0085
R3582 X2.n457 X2.n300 0.0085
R3583 X2.n746 X2.n9 0.0085
R3584 X2.n1141 X2.n142 0.00809524
R3585 X2.n730 X2.n539 0.00778095
R3586 X2.n1212 X2.n109 0.00763514
R3587 X2.n1299 X2.n67 0.00763514
R3588 X2.n466 X2.n350 0.00763514
R3589 X2.n537 X2.n13 0.00763514
R3590 X2.n708 X2.n23 0.00741892
R3591 X2.n624 X2.n623 0.00741892
R3592 X2.n846 X2.n262 0.00741892
R3593 X2.n1050 X2.n169 0.00741892
R3594 X2.n1187 X2.n119 0.00741892
R3595 X2.n1277 X2.n1276 0.00741892
R3596 X2.n450 X2.n356 0.00741892
R3597 X2.n525 X2.n8 0.00741892
R3598 X2.n750 X2.n523 0.00725714
R3599 X2.n730 X2.n729 0.00707381
R3600 X2.n722 X2.n18 0.00698649
R3601 X2.n607 X2.n605 0.00698649
R3602 X2.n813 X2.n281 0.00698649
R3603 X2.n1098 X2.n1097 0.00698649
R3604 X2.n391 X2.n370 0.00696162
R3605 X2.n602 X2.n600 0.00691667
R3606 X2.n677 X2.n676 0.00666216
R3607 X2.n655 X2.n38 0.00666216
R3608 X2.n237 X2.n224 0.00666216
R3609 X2.n977 X2.n976 0.00666216
R3610 X2.n1214 X2.n107 0.00655405
R3611 X2.n1312 X2.n62 0.00655405
R3612 X2.n473 X2.n305 0.00655405
R3613 X2.n733 X2.n14 0.00655405
R3614 X2.n1182 X2.n1181 0.00633784
R3615 X2.n1282 X2.n1281 0.00633784
R3616 X2.n445 X2.n297 0.00633784
R3617 X2.n518 X2.n517 0.00633784
R3618 X2.n568 X2.n29 0.00590541
R3619 X2.n644 X2.n40 0.00590541
R3620 X2.n243 X2.n242 0.00590541
R3621 X2.n198 X2.n192 0.00590541
R3622 X2.n490 X2.n339 0.00588776
R3623 X2.n401 X2.n370 0.00588776
R3624 X2.n1220 X2.n1219 0.00547297
R3625 X2.n1313 X2.n55 0.00547297
R3626 X2.n475 X2.n306 0.00547297
R3627 X2.n542 X2.n15 0.00547297
R3628 X2.n129 X2.n128 0.00525676
R3629 X2.n1268 X2.n1267 0.00525676
R3630 X2.n438 X2.n296 0.00525676
R3631 X2.n757 X2.n756 0.00525676
R3632 X2.n697 X2.n25 0.00514865
R3633 X2.n591 X2.n44 0.00514865
R3634 X2.n871 X2.n254 0.00514865
R3635 X2.n1033 X2.n177 0.00514865
R3636 X2.n1318 X2.n59 0.00440238
R3637 X2.n663 X2.n35 0.00439189
R3638 X2.n217 X2.n212 0.00439189
R3639 X2.n1117 X2.n150 0.00439189
R3640 X2.n1228 X2.n96 0.00439189
R3641 X2.n393 X2.n286 0.00439189
R3642 X2.n484 X2.n307 0.00439189
R3643 X2.n724 X2.n723 0.00425921
R3644 X2.n720 X2.n719 0.00425921
R3645 X2.n706 X2.n703 0.00425921
R3646 X2.n561 X2.n553 0.00425921
R3647 X2.n692 X2.n691 0.00425921
R3648 X2.n569 X2.n565 0.00425921
R3649 X2.n685 X2.n682 0.00425921
R3650 X2.n680 X2.n570 0.00425921
R3651 X2.n665 X2.n662 0.00425921
R3652 X2.n653 X2.n650 0.00425921
R3653 X2.n584 X2.n578 0.00425921
R3654 X2.n645 X2.n585 0.00425921
R3655 X2.n640 X2.n639 0.00425921
R3656 X2.n632 X2.n629 0.00425921
R3657 X2.n627 X2.n593 0.00425921
R3658 X2.n610 X2.n609 0.00425921
R3659 X2.n606 X2.n56 0.00425921
R3660 X2.n144 X2.n141 0.00425921
R3661 X2.n1148 X2.n1147 0.00425921
R3662 X2.n1144 X2.n132 0.00425921
R3663 X2.n1161 X2.n134 0.00425921
R3664 X2.n1186 X2.n1184 0.00425921
R3665 X2.n1191 X2.n118 0.00425921
R3666 X2.n1202 X2.n115 0.00425921
R3667 X2.n1196 X2.n116 0.00425921
R3668 X2.n1222 X2.n98 0.00425921
R3669 X2.n1238 X2.n91 0.00425921
R3670 X2.n1249 X2.n88 0.00425921
R3671 X2.n1243 X2.n89 0.00425921
R3672 X2.n1244 X2.n81 0.00425921
R3673 X2.n1279 X2.n1278 0.00425921
R3674 X2.n1274 X2.n70 0.00425921
R3675 X2.n1293 X2.n68 0.00425921
R3676 X2.n1304 X2.n1298 0.00425921
R3677 X2.n453 X2.n452 0.00425921
R3678 X2.n459 X2.n456 0.00425921
R3679 X2.n528 X2.n527 0.00425921
R3680 X2.n748 X2.n745 0.00425921
R3681 X2.n740 X2.n533 0.00424524
R3682 X2.n719 X2.n548 0.0042371
R3683 X2.n715 X2.n714 0.0042371
R3684 X2.n711 X2.n710 0.0042371
R3685 X2.n707 X2.n706 0.0042371
R3686 X2.n698 X2.n562 0.0042371
R3687 X2.n693 X2.n692 0.0042371
R3688 X2.n675 X2.n570 0.0042371
R3689 X2.n574 X2.n572 0.0042371
R3690 X2.n670 X2.n666 0.0042371
R3691 X2.n666 X2.n665 0.0042371
R3692 X2.n662 X2.n661 0.0042371
R3693 X2.n658 X2.n657 0.0042371
R3694 X2.n654 X2.n653 0.0042371
R3695 X2.n639 X2.n638 0.0042371
R3696 X2.n592 X2.n588 0.0042371
R3697 X2.n622 X2.n593 0.0042371
R3698 X2.n597 X2.n595 0.0042371
R3699 X2.n617 X2.n614 0.0042371
R3700 X2.n611 X2.n610 0.0042371
R3701 X2.n1120 X2.n143 0.0042371
R3702 X2.n1139 X2.n144 0.0042371
R3703 X2.n134 X2.n133 0.0042371
R3704 X2.n1171 X2.n1170 0.0042371
R3705 X2.n1165 X2.n130 0.0042371
R3706 X2.n1184 X2.n120 0.0042371
R3707 X2.n1197 X2.n1196 0.0042371
R3708 X2.n1215 X2.n108 0.0042371
R3709 X2.n1217 X2.n106 0.0042371
R3710 X2.n1222 X2.n106 0.0042371
R3711 X2.n1226 X2.n98 0.0042371
R3712 X2.n104 X2.n103 0.0042371
R3713 X2.n99 X2.n91 0.0042371
R3714 X2.n1262 X2.n81 0.0042371
R3715 X2.n1264 X2.n79 0.0042371
R3716 X2.n1269 X2.n77 0.0042371
R3717 X2.n1280 X2.n1279 0.0042371
R3718 X2.n1304 X2.n1303 0.0042371
R3719 X2.n1301 X2.n61 0.0042371
R3720 X2.n1315 X2.n57 0.0042371
R3721 X2.n1319 X2.n57 0.0042371
R3722 X2.n411 X2.n404 0.0042371
R3723 X2.n436 X2.n433 0.0042371
R3724 X2.n439 X2.n358 0.0042371
R3725 X2.n477 X2.n347 0.0042371
R3726 X2.n497 X2.n344 0.0042371
R3727 X2.n325 X2.n323 0.0042371
R3728 X2.n755 X2.n754 0.0042371
R3729 X2.n735 X2.n732 0.0042371
R3730 X2.n543 X2.n540 0.0042371
R3731 X2.n1126 X2.n1125 0.00423273
R3732 X2.n481 X2.n347 0.00423268
R3733 X2.n1114 X2.n1113 0.00422178
R3734 X2.n376 X2.n373 0.00422178
R3735 X2.n532 X2.n523 0.00421905
R3736 X2.n1173 X2.n1172 0.00417568
R3737 X2.n1265 X2.n80 0.00417568
R3738 X2.n434 X2.n295 0.00417568
R3739 X2.n324 X2.n316 0.00417568
R3740 X2.n715 X2.n549 0.00410442
R3741 X2.n614 X2.n598 0.00410442
R3742 X2.n712 X2.n551 0.00406757
R3743 X2.n615 X2.n48 0.00406757
R3744 X2.n837 X2.n266 0.00406757
R3745 X2.n1090 X2.n1089 0.00406757
R3746 X2.n474 X2.n349 0.00402269
R3747 X2.n368 X2.n364 0.00398793
R3748 X2.n337 X2.n333 0.00398793
R3749 X2.n1148 X2.n1143 0.00397174
R3750 X2.n1202 X2.n1201 0.00397174
R3751 X2.n1239 X2.n88 0.00397174
R3752 X2.n1297 X2.n68 0.00397174
R3753 X2.n682 X2.n681 0.00394963
R3754 X2.n649 X2.n578 0.00394963
R3755 X2.n403 X2.n402 0.00394626
R3756 X2.n491 X2.n340 0.00394626
R3757 X2.n395 X2.n394 0.00393696
R3758 X2.n486 X2.n485 0.00393696
R3759 X2.n419 X2.n418 0.00390294
R3760 X2.n506 X2.n502 0.00390294
R3761 X2.n464 X2.n351 0.00389381
R3762 X2.n428 X2.n427 0.00385851
R3763 X2.n448 X2.n447 0.00385851
R3764 X2.n332 X2.n331 0.00385851
R3765 X2.n521 X2.n520 0.00385851
R3766 X2.n428 X2.n360 0.00380768
R3767 X2.n331 X2.n322 0.00380768
R3768 X2.n447 X2.n357 0.00380053
R3769 X2.n520 X2.n321 0.00380053
R3770 X2.n702 X2.n553 0.00379484
R3771 X2.n629 X2.n628 0.00379484
R3772 X2.n1127 X2.n153 0.00379484
R3773 X2.n727 X2.n544 0.00377273
R3774 X2.n404 X2.n366 0.0037725
R3775 X2.n464 X2.n463 0.0037725
R3776 X2.n344 X2.n335 0.0037725
R3777 X2.n739 X2.n738 0.00374762
R3778 X2.n1171 X2.n127 0.0037285
R3779 X2.n1264 X2.n1263 0.0037285
R3780 X2.n1166 X2.n1165 0.00370639
R3781 X2.n1273 X2.n77 0.00370639
R3782 X2.n737 X2.n539 0.00369524
R3783 X2.n564 X2.n562 0.00366216
R3784 X2.n636 X2.n588 0.00366216
R3785 X2.n742 X2.n741 0.00366216
R3786 X2.n531 X2.n529 0.00364005
R3787 X2.n718 X2.n19 0.00363514
R3788 X2.n599 X2.n50 0.00363514
R3789 X2.n811 X2.n274 0.00363514
R3790 X2.n1096 X2.n159 0.00363514
R3791 X2.n1124 X2.n1123 0.00359048
R3792 X2.n456 X2.n353 0.00358532
R3793 X2.n482 X2.n346 0.00358218
R3794 X2.n377 X2.n376 0.00357902
R3795 X2.n1113 X2.n154 0.00357902
R3796 X2.n369 X2.n368 0.00357098
R3797 X2.n338 X2.n337 0.00357098
R3798 X2.n689 X2.n565 0.00348526
R3799 X2.n587 X2.n585 0.00348526
R3800 X2.n433 X2.n432 0.003457
R3801 X2.n326 X2.n325 0.003457
R3802 X2.n443 X2.n358 0.00344926
R3803 X2.n754 X2.n753 0.00344926
R3804 X2.n1162 X2.n132 0.00344103
R3805 X2.n1185 X2.n118 0.00344103
R3806 X2.n1245 X2.n1243 0.00344103
R3807 X2.n1275 X2.n1274 0.00344103
R3808 X2.n449 X2.n355 0.00343273
R3809 X2.n524 X2.n522 0.00343273
R3810 X2.n363 X2.n362 0.00341839
R3811 X2.n504 X2.n327 0.00341839
R3812 X2.n513 X2.n334 0.00341837
R3813 X2.n425 X2.n365 0.00341837
R3814 X2.n1122 X2.n142 0.00335476
R3815 X2.n710 X2.n552 0.00335258
R3816 X2.n621 X2.n595 0.00335258
R3817 X2.n418 X2.n363 0.0033136
R3818 X2.n506 X2.n327 0.0033136
R3819 X2.n667 X2.n33 0.00331081
R3820 X2.n659 X2.n576 0.00331081
R3821 X2.n933 X2.n931 0.00331081
R3822 X2.n962 X2.n961 0.00331081
R3823 X2.n1134 X2.n145 0.00331081
R3824 X2.n101 X2.n97 0.00331081
R3825 X2.n396 X2.n287 0.00331081
R3826 X2.n494 X2.n493 0.00331081
R3827 X2.n444 X2.n443 0.00330444
R3828 X2.n753 X2.n320 0.00330444
R3829 X2.n452 X2.n355 0.0032992
R3830 X2.n527 X2.n522 0.0032992
R3831 X2.n432 X2.n431 0.00329663
R3832 X2.n328 X2.n326 0.00329663
R3833 X2.n538 X2.n535 0.00324201
R3834 X2.n674 X2.n572 0.00319779
R3835 X2.n657 X2.n577 0.00319779
R3836 X2.n1198 X2.n108 0.00319779
R3837 X2.n1302 X2.n1301 0.00319779
R3838 X2.n736 X2.n735 0.00319779
R3839 X2.n1140 X2.n143 0.00317568
R3840 X2.n103 X2.n100 0.00317568
R3841 X2.n412 X2.n403 0.00317568
R3842 X2.n498 X2.n340 0.00317568
R3843 X2.n406 X2.n369 0.00316007
R3844 X2.n341 X2.n338 0.00316007
R3845 X2.n353 X2.n352 0.00314581
R3846 X2.n1119 X2.n1116 0.00310934
R3847 X2.n1159 X2.n1158 0.00309459
R3848 X2.n1260 X2.n1259 0.00309459
R3849 X2.n429 X2.n361 0.00309459
R3850 X2.n330 X2.n315 0.00309459
R3851 X2.n723 X2.n547 0.003043
R3852 X2.n606 X2.n604 0.003043
R3853 X2.n842 X2.n840 0.0029881
R3854 X2.n875 X2.n252 0.0029881
R3855 X2.n898 X2.n890 0.0029881
R3856 X2.n1014 X2.n1013 0.0029881
R3857 X2.n406 X2.n366 0.00298054
R3858 X2.n463 X2.n352 0.00298054
R3859 X2.n341 X2.n335 0.00298054
R3860 X2.n1029 X2.n180 0.0029619
R3861 X2.n1061 X2.n1060 0.0029619
R3862 X2.n444 X2.n357 0.00293083
R3863 X2.n321 X2.n320 0.00293083
R3864 X2.n431 X2.n360 0.0029237
R3865 X2.n328 X2.n322 0.0029237
R3866 X2.n671 X2.n574 0.00291032
R3867 X2.n658 X2.n575 0.00291032
R3868 X2.n1121 X2.n1120 0.00291032
R3869 X2.n1216 X2.n1215 0.00291032
R3870 X2.n1225 X2.n104 0.00291032
R3871 X2.n1316 X2.n61 0.00291032
R3872 X2.n478 X2.n474 0.00291032
R3873 X2.n732 X2.n731 0.00291032
R3874 X2.n427 X2.n362 0.00289527
R3875 X2.n449 X2.n448 0.00289527
R3876 X2.n504 X2.n332 0.00289527
R3877 X2.n524 X2.n521 0.00289527
R3878 X2.n378 X2.n377 0.00287188
R3879 X2.n1111 X2.n154 0.00284569
R3880 X2.n467 X2.n351 0.00283826
R3881 X2.n600 X2.n59 0.00283095
R3882 X2.n398 X2.n395 0.00279542
R3883 X2.n487 X2.n486 0.00279542
R3884 X2.n415 X2.n364 0.00276679
R3885 X2.n501 X2.n333 0.00276679
R3886 X2.n711 X2.n550 0.00275553
R3887 X2.n618 X2.n597 0.00275553
R3888 X2.n724 X2.n546 0.00273342
R3889 X2.n1319 X2.n56 0.00273342
R3890 X2.n386 X2.n378 0.00272619
R3891 X2.n386 X2.n385 0.00272619
R3892 X2.n816 X2.n279 0.00272619
R3893 X2.n818 X2.n817 0.00272619
R3894 X2.n826 X2.n825 0.00272619
R3895 X2.n834 X2.n268 0.00272619
R3896 X2.n839 X2.n268 0.00272619
R3897 X2.n841 X2.n264 0.00272619
R3898 X2.n849 X2.n264 0.00272619
R3899 X2.n851 X2.n260 0.00272619
R3900 X2.n859 X2.n260 0.00272619
R3901 X2.n867 X2.n256 0.00272619
R3902 X2.n868 X2.n867 0.00272619
R3903 X2.n877 X2.n876 0.00272619
R3904 X2.n877 X2.n248 0.00272619
R3905 X2.n885 X2.n246 0.00272619
R3906 X2.n889 X2.n246 0.00272619
R3907 X2.n897 X2.n896 0.00272619
R3908 X2.n892 X2.n891 0.00272619
R3909 X2.n915 X2.n229 0.00272619
R3910 X2.n925 X2.n924 0.00272619
R3911 X2.n928 X2.n925 0.00272619
R3912 X2.n936 X2.n222 0.00272619
R3913 X2.n937 X2.n936 0.00272619
R3914 X2.n938 X2.n937 0.00272619
R3915 X2.n952 X2.n951 0.00272619
R3916 X2.n966 X2.n210 0.00272619
R3917 X2.n967 X2.n966 0.00272619
R3918 X2.n973 X2.n972 0.00272619
R3919 X2.n974 X2.n973 0.00272619
R3920 X2.n974 X2.n204 0.00272619
R3921 X2.n983 X2.n202 0.00272619
R3922 X2.n987 X2.n202 0.00272619
R3923 X2.n993 X2.n992 0.00272619
R3924 X2.n992 X2.n989 0.00272619
R3925 X2.n1019 X2.n188 0.00272619
R3926 X2.n1028 X2.n1027 0.00272619
R3927 X2.n1036 X2.n1035 0.00272619
R3928 X2.n1038 X2.n1037 0.00272619
R3929 X2.n1047 X2.n1046 0.00272619
R3930 X2.n1056 X2.n167 0.00272619
R3931 X2.n1060 X2.n167 0.00272619
R3932 X2.n1087 X2.n1086 0.00272619
R3933 X2.n1086 X2.n1085 0.00272619
R3934 X2.n1085 X2.n1062 0.00272619
R3935 X2.n1076 X2.n1064 0.00272619
R3936 X2.n1076 X2.n1075 0.00272619
R3937 X2.n1069 X2.n157 0.00272619
R3938 X2.n1102 X2.n157 0.00272619
R3939 X2.n1109 X2.n1108 0.00272619
R3940 X2.n1111 X2.n1110 0.00272619
R3941 X2.n385 X2.n384 0.0027
R3942 X2.n817 X2.n816 0.0027
R3943 X2.n826 X2.n824 0.0027
R3944 X2.n834 X2.n833 0.0027
R3945 X2.n842 X2.n841 0.0027
R3946 X2.n869 X2.n868 0.0027
R3947 X2.n896 X2.n891 0.0027
R3948 X2.n915 X2.n914 0.0027
R3949 X2.n924 X2.n227 0.0027
R3950 X2.n952 X2.n944 0.0027
R3951 X2.n945 X2.n210 0.0027
R3952 X2.n989 X2.n190 0.0027
R3953 X2.n1015 X2.n188 0.0027
R3954 X2.n1027 X2.n184 0.0027
R3955 X2.n1038 X2.n1036 0.0027
R3956 X2.n1047 X2.n1045 0.0027
R3957 X2.n1056 X2.n1055 0.0027
R3958 X2.n1103 X2.n1102 0.0027
R3959 X2.n1110 X2.n1109 0.0027
R3960 X2.n869 X2.n252 0.00264762
R3961 X2.n1035 X2.n180 0.00264762
R3962 X2.n1145 X2.n1144 0.00264496
R3963 X2.n1248 X2.n89 0.00264496
R3964 X2.n1192 X2.n1191 0.00262285
R3965 X2.n1294 X2.n70 0.00262285
R3966 X2.n460 X2.n453 0.00262285
R3967 X2.n749 X2.n528 0.00262285
R3968 X2.n890 X2.n889 0.00262143
R3969 X2.n1015 X2.n1014 0.00262143
R3970 X2.n686 X2.n569 0.00260074
R3971 X2.n646 X2.n645 0.00260074
R3972 X2.n844 X2.n267 0.00257862
R3973 X2.n1059 X2.n165 0.00257862
R3974 X2.n1013 X2.n190 0.00256905
R3975 X2.n690 X2.n28 0.00255405
R3976 X2.n642 X2.n641 0.00255405
R3977 X2.n902 X2.n241 0.00255405
R3978 X2.n1009 X2.n186 0.00255405
R3979 X2.n898 X2.n897 0.00254286
R3980 X2.n1029 X2.n1028 0.00254286
R3981 X2.n900 X2.n899 0.0025344
R3982 X2.n876 X2.n875 0.00251667
R3983 X2.n1012 X2.n1011 0.00251228
R3984 X2.n482 X2.n481 0.00249519
R3985 X2.n390 X2.n389 0.0024936
R3986 X2.n840 X2.n839 0.00246429
R3987 X2.n1087 X2.n1061 0.00246429
R3988 X2.n699 X2.n698 0.00244595
R3989 X2.n633 X2.n592 0.00244595
R3990 X2.n860 X2.n859 0.0024381
R3991 X2.n1045 X2.n1044 0.0024381
R3992 X2.n873 X2.n253 0.00242383
R3993 X2.n1031 X2.n181 0.00242383
R3994 X2.n740 X2.n739 0.00238571
R3995 X2.n1125 X2.n1124 0.00238571
R3996 X2.n823 X2.n277 0.00238571
R3997 X2.n832 X2.n272 0.00238571
R3998 X2.n852 X2.n850 0.00238571
R3999 X2.n861 X2.n860 0.00238571
R4000 X2.n884 X2.n883 0.00238571
R4001 X2.n913 X2.n232 0.00238571
R4002 X2.n920 X2.n919 0.00238571
R4003 X2.n943 X2.n220 0.00238571
R4004 X2.n950 X2.n946 0.00238571
R4005 X2.n968 X2.n967 0.00238571
R4006 X2.n982 X2.n981 0.00238571
R4007 X2.n994 X2.n988 0.00238571
R4008 X2.n1021 X2.n1020 0.00238571
R4009 X2.n1044 X2.n175 0.00238571
R4010 X2.n1054 X2.n170 0.00238571
R4011 X2.n1081 X2.n1080 0.00238571
R4012 X2.n1074 X2.n1070 0.00238571
R4013 X2.n815 X2.n814 0.00237961
R4014 X2.n819 X2.n278 0.00237961
R4015 X2.n827 X2.n276 0.00237961
R4016 X2.n835 X2.n269 0.00237961
R4017 X2.n838 X2.n269 0.00237961
R4018 X2.n847 X2.n265 0.00237961
R4019 X2.n848 X2.n847 0.00237961
R4020 X2.n857 X2.n261 0.00237961
R4021 X2.n858 X2.n857 0.00237961
R4022 X2.n866 X2.n257 0.00237961
R4023 X2.n866 X2.n255 0.00237961
R4024 X2.n878 X2.n251 0.00237961
R4025 X2.n878 X2.n249 0.00237961
R4026 X2.n887 X2.n886 0.00237961
R4027 X2.n888 X2.n887 0.00237961
R4028 X2.n895 X2.n245 0.00237961
R4029 X2.n894 X2.n893 0.00237961
R4030 X2.n917 X2.n916 0.00237961
R4031 X2.n923 X2.n225 0.00237961
R4032 X2.n929 X2.n225 0.00237961
R4033 X2.n935 X2.n934 0.00237961
R4034 X2.n935 X2.n221 0.00237961
R4035 X2.n939 X2.n221 0.00237961
R4036 X2.n953 X2.n219 0.00237961
R4037 X2.n965 X2.n964 0.00237961
R4038 X2.n965 X2.n209 0.00237961
R4039 X2.n971 X2.n207 0.00237961
R4040 X2.n975 X2.n207 0.00237961
R4041 X2.n975 X2.n205 0.00237961
R4042 X2.n985 X2.n984 0.00237961
R4043 X2.n986 X2.n985 0.00237961
R4044 X2.n991 X2.n201 0.00237961
R4045 X2.n991 X2.n990 0.00237961
R4046 X2.n1018 X2.n1017 0.00237961
R4047 X2.n1026 X2.n183 0.00237961
R4048 X2.n1034 X2.n178 0.00237961
R4049 X2.n1039 X2.n179 0.00237961
R4050 X2.n1048 X2.n174 0.00237961
R4051 X2.n1058 X2.n1057 0.00237961
R4052 X2.n1059 X2.n1058 0.00237961
R4053 X2.n1088 X2.n166 0.00237961
R4054 X2.n1084 X2.n166 0.00237961
R4055 X2.n1084 X2.n1083 0.00237961
R4056 X2.n1078 X2.n1077 0.00237961
R4057 X2.n1077 X2.n1068 0.00237961
R4058 X2.n1100 X2.n158 0.00237961
R4059 X2.n1101 X2.n1100 0.00237961
R4060 X2.n1107 X2.n151 0.00237961
R4061 X2.n1170 X2.n1169 0.00237961
R4062 X2.n1169 X2.n130 0.00237961
R4063 X2.n1270 X2.n79 0.00237961
R4064 X2.n1270 X2.n1269 0.00237961
R4065 X2.n388 X2.n372 0.00237961
R4066 X2.n400 X2.n371 0.00237961
R4067 X2.n440 X2.n436 0.00237961
R4068 X2.n440 X2.n439 0.00237961
R4069 X2.n471 X2.n470 0.00237961
R4070 X2.n492 X2.n489 0.00237961
R4071 X2.n323 X2.n319 0.00237961
R4072 X2.n755 X2.n319 0.00237961
R4073 X2.n914 X2.n913 0.00235952
R4074 X2.n926 X2.n222 0.00235952
R4075 X2.n383 X2.n374 0.00235749
R4076 X2.n815 X2.n278 0.00235749
R4077 X2.n827 X2.n275 0.00235749
R4078 X2.n835 X2.n271 0.00235749
R4079 X2.n843 X2.n265 0.00235749
R4080 X2.n870 X2.n255 0.00235749
R4081 X2.n895 X2.n894 0.00235749
R4082 X2.n916 X2.n230 0.00235749
R4083 X2.n923 X2.n922 0.00235749
R4084 X2.n953 X2.n218 0.00235749
R4085 X2.n964 X2.n211 0.00235749
R4086 X2.n990 X2.n191 0.00235749
R4087 X2.n1017 X2.n1016 0.00235749
R4088 X2.n1026 X2.n185 0.00235749
R4089 X2.n1039 X2.n178 0.00235749
R4090 X2.n1048 X2.n173 0.00235749
R4091 X2.n1057 X2.n168 0.00235749
R4092 X2.n1101 X2.n156 0.00235749
R4093 X2.n423 X2.n422 0.00235749
R4094 X2.n511 X2.n510 0.00235749
R4095 X2.n988 X2.n987 0.00233333
R4096 X2.n870 X2.n253 0.00231327
R4097 X2.n1034 X2.n181 0.00231327
R4098 X2.n384 X2.n380 0.00230714
R4099 X2.n1104 X2.n1103 0.00230714
R4100 X2.n1108 X2.n155 0.00230714
R4101 X2.n699 X2.n561 0.00229115
R4102 X2.n633 X2.n632 0.00229115
R4103 X2.n888 X2.n244 0.00229115
R4104 X2.n1016 X2.n189 0.00229115
R4105 X2.n379 X2.n279 0.00228095
R4106 X2.n825 X2.n272 0.00228095
R4107 X2.n1080 X2.n1064 0.00225476
R4108 X2.n1012 X2.n191 0.00224693
R4109 X2.n1138 X2.n1137 0.00222973
R4110 X2.n1234 X2.n92 0.00222973
R4111 X2.n410 X2.n409 0.00222973
R4112 X2.n496 X2.n310 0.00222973
R4113 X2.n899 X2.n245 0.00222482
R4114 X2.n1030 X2.n183 0.00222482
R4115 X2.n874 X2.n251 0.0022027
R4116 X2.n928 X2.n927 0.00220238
R4117 X2.n972 X2.n208 0.00220238
R4118 X2.n944 X2.n943 0.00217619
R4119 X2.n951 X2.n950 0.00217619
R4120 X2.n485 X2.n346 0.00217613
R4121 X2.n838 X2.n267 0.00215848
R4122 X2.n1088 X2.n165 0.00215848
R4123 X2.n686 X2.n685 0.00213636
R4124 X2.n646 X2.n584 0.00213636
R4125 X2.n858 X2.n259 0.00213636
R4126 X2.n1043 X2.n173 0.00213636
R4127 X2.n1192 X2.n115 0.00211425
R4128 X2.n1294 X2.n1293 0.00211425
R4129 X2.n460 X2.n459 0.00211425
R4130 X2.n749 X2.n748 0.00211425
R4131 X2.n1123 X2.n1122 0.00209762
R4132 X2.n824 X2.n823 0.00209762
R4133 X2.n969 X2.n209 0.00209214
R4134 X2.n1147 X2.n1145 0.00209214
R4135 X2.n1249 X2.n1248 0.00209214
R4136 X2.n424 X2.n415 0.00209214
R4137 X2.n512 X2.n501 0.00209214
R4138 X2.n1075 X2.n1074 0.00207143
R4139 X2.n912 X2.n230 0.00207002
R4140 X2.n934 X2.n223 0.00207002
R4141 X2.n986 X2.n200 0.00204791
R4142 X2.n383 X2.n382 0.0020258
R4143 X2.n1105 X2.n156 0.0020258
R4144 X2.n1107 X2.n1106 0.0020258
R4145 X2.n919 X2.n229 0.00201905
R4146 X2.n1157 X2.n1156 0.00201351
R4147 X2.n1242 X2.n1241 0.00201351
R4148 X2.n417 X2.n292 0.00201351
R4149 X2.n508 X2.n507 0.00201351
R4150 X2.n714 X2.n550 0.00200369
R4151 X2.n618 X2.n617 0.00200369
R4152 X2.n814 X2.n280 0.00200369
R4153 X2.n276 X2.n273 0.00200369
R4154 X2.n1126 X2.n1114 0.00200107
R4155 X2.n389 X2.n373 0.00200107
R4156 X2.n391 X2.n390 0.00200107
R4157 X2.n983 X2.n982 0.00199286
R4158 X2.n1079 X2.n1078 0.00198157
R4159 X2.n929 X2.n226 0.00193735
R4160 X2.n971 X2.n970 0.00193735
R4161 X2.n942 X2.n218 0.00191523
R4162 X2.n949 X2.n219 0.00191523
R4163 X2.n1127 X2.n152 0.00191523
R4164 X2.n1319 X2.n58 0.00191523
R4165 X2.n388 X2.n387 0.00191523
R4166 X2.n392 X2.n372 0.00191523
R4167 X2.n852 X2.n851 0.00191429
R4168 X2.n1046 X2.n170 0.00191429
R4169 X2.n863 X2.n862 0.00187101
R4170 X2.n422 X2.n419 0.00185493
R4171 X2.n510 X2.n502 0.00185493
R4172 X2.n671 X2.n670 0.00184889
R4173 X2.n661 X2.n575 0.00184889
R4174 X2.n822 X2.n275 0.00184889
R4175 X2.n1042 X2.n176 0.00184889
R4176 X2.n1121 X2.n1119 0.00184889
R4177 X2.n1217 X2.n1216 0.00184889
R4178 X2.n1226 X2.n1225 0.00184889
R4179 X2.n1316 X2.n1315 0.00184889
R4180 X2.n399 X2.n398 0.00184889
R4181 X2.n478 X2.n477 0.00184889
R4182 X2.n488 X2.n487 0.00184889
R4183 X2.n731 X2.n540 0.00184889
R4184 X2.n1021 X2.n184 0.00183571
R4185 X2.n1073 X2.n1068 0.00182678
R4186 X2.n883 X2.n248 0.00180952
R4187 X2.n695 X2.n694 0.0017973
R4188 X2.n637 X2.n43 0.0017973
R4189 X2.n879 X2.n250 0.0017973
R4190 X2.n1025 X2.n182 0.0017973
R4191 X2.n402 X2.n371 0.0017897
R4192 X2.n492 X2.n491 0.0017897
R4193 X2.n911 X2.n233 0.00178256
R4194 X2.n918 X2.n917 0.00178256
R4195 X2.n996 X2.n995 0.00178256
R4196 X2.n984 X2.n203 0.00176044
R4197 X2.n738 X2.n737 0.00175714
R4198 X2.n885 X2.n884 0.00173095
R4199 X2.n1020 X2.n1019 0.00173095
R4200 X2.n831 X2.n830 0.00171622
R4201 X2.n471 X2.n349 0.00171347
R4202 X2.n720 X2.n547 0.0016941
R4203 X2.n609 X2.n604 0.0016941
R4204 X2.n853 X2.n261 0.0016941
R4205 X2.n174 X2.n171 0.0016941
R4206 X2.n1082 X2.n1063 0.0016941
R4207 X2.n1055 X2.n1054 0.00165238
R4208 X2.n941 X2.n940 0.00162776
R4209 X2.n948 X2.n947 0.00162776
R4210 X2.n1022 X2.n185 0.00162776
R4211 X2.n1116 X2.n1115 0.00162776
R4212 X2.n850 X2.n849 0.00162619
R4213 X2.n882 X2.n249 0.00160565
R4214 X2.n1140 X2.n1139 0.00158354
R4215 X2.n100 X2.n99 0.00158354
R4216 X2.n412 X2.n411 0.00158354
R4217 X2.n498 X2.n497 0.00158354
R4218 X2.n675 X2.n674 0.00156143
R4219 X2.n654 X2.n577 0.00156143
R4220 X2.n821 X2.n820 0.00156143
R4221 X2.n1072 X2.n1071 0.00156143
R4222 X2.n1198 X2.n1197 0.00156143
R4223 X2.n1303 X2.n1302 0.00156143
R4224 X2.n468 X2.n467 0.00156143
R4225 X2.n736 X2.n538 0.00156143
R4226 X2.n920 X2.n227 0.00154762
R4227 X2.n981 X2.n204 0.00154762
R4228 X2.n886 X2.n247 0.00153931
R4229 X2.n1018 X2.n187 0.00153931
R4230 X2.n921 X2.n228 0.00149509
R4231 X2.n535 X2.n534 0.00149509
R4232 X2.n980 X2.n979 0.00147297
R4233 X2.n1053 X2.n168 0.00147297
R4234 X2.n818 X2.n277 0.00146905
R4235 X2.n1070 X2.n1069 0.00146905
R4236 X2.n848 X2.n263 0.00145086
R4237 X2.n707 X2.n552 0.00140663
R4238 X2.n622 X2.n621 0.00140663
R4239 X2.n854 X2.n263 0.00140663
R4240 X2.n1053 X2.n1052 0.00140663
R4241 X2.n946 X2.n945 0.00139048
R4242 X2.n922 X2.n921 0.00138452
R4243 X2.n980 X2.n205 0.00138452
R4244 X2.n380 X2.n379 0.00136429
R4245 X2.n927 X2.n926 0.00136429
R4246 X2.n938 X2.n220 0.00136429
R4247 X2.n881 X2.n247 0.00134029
R4248 X2.n1023 X2.n187 0.00134029
R4249 X2.n968 X2.n208 0.00133809
R4250 X2.n1104 X2.n155 0.00133809
R4251 X2.n820 X2.n819 0.00131818
R4252 X2.n1071 X2.n158 0.00131818
R4253 X2.n470 X2.n468 0.00131818
R4254 X2.n1162 X2.n1161 0.00129607
R4255 X2.n1186 X2.n1185 0.00129607
R4256 X2.n1245 X2.n1244 0.00129607
R4257 X2.n1278 X2.n1275 0.00129607
R4258 X2.n833 X2.n832 0.00128571
R4259 X2.n1081 X2.n1062 0.00128571
R4260 X2.n691 X2.n689 0.00125184
R4261 X2.n640 X2.n587 0.00125184
R4262 X2.n882 X2.n881 0.00125184
R4263 X2.n947 X2.n211 0.00125184
R4264 X2.n1023 X2.n1022 0.00125184
R4265 X2.n382 X2.n280 0.00122973
R4266 X2.n226 X2.n223 0.00122973
R4267 X2.n940 X2.n939 0.00122973
R4268 X2.n970 X2.n969 0.00120762
R4269 X2.n1106 X2.n1105 0.00120762
R4270 X2.n892 X2.n232 0.00120714
R4271 X2.n994 X2.n993 0.00120714
R4272 X2.n854 X2.n853 0.0011855
R4273 X2.n1052 X2.n171 0.0011855
R4274 X2.n831 X2.n271 0.00116339
R4275 X2.n1083 X2.n1082 0.00116339
R4276 X2.n1150 X2.n139 0.00114865
R4277 X2.n1237 X2.n1236 0.00114865
R4278 X2.n407 X2.n290 0.00114865
R4279 X2.n342 X2.n311 0.00114865
R4280 X2.n1037 X2.n175 0.00112857
R4281 X2.n979 X2.n203 0.00111916
R4282 X2.n861 X2.n256 0.00110238
R4283 X2.n693 X2.n564 0.00109705
R4284 X2.n638 X2.n636 0.00109705
R4285 X2.n893 X2.n233 0.00109705
R4286 X2.n918 X2.n228 0.00109705
R4287 X2.n995 X2.n201 0.00109705
R4288 X2.n741 X2.n534 0.00109705
R4289 X2.n1166 X2.n120 0.00105283
R4290 X2.n1280 X2.n1273 0.00105283
R4291 X2.n601 X2.n58 0.00105283
R4292 X2.n668 X2.n34 0.00104054
R4293 X2.n955 X2.n216 0.00104054
R4294 X2.n822 X2.n821 0.00103071
R4295 X2.n179 X2.n176 0.00103071
R4296 X2.n1073 X2.n1072 0.00103071
R4297 X2.n1112 X2.n152 0.00103071
R4298 X2.n133 X2.n127 0.00103071
R4299 X2.n1263 X2.n1262 0.00103071
R4300 X2.n387 X2.n375 0.00103071
R4301 X2.n400 X2.n399 0.00103071
R4302 X2.n489 X2.n488 0.00103071
R4303 X2.n862 X2.n257 0.0010086
R4304 X2.n942 X2.n941 0.000964373
R4305 X2.n949 X2.n948 0.000964373
R4306 X2.n1115 X2.n153 0.000964373
R4307 X2.n394 X2.n392 0.000964373
R4308 X2.n544 X2.n543 0.000964373
R4309 X2.n703 X2.n702 0.00094226
R4310 X2.n628 X2.n627 0.00094226
R4311 X2.n1146 X2.n140 0.000932432
R4312 X2.n1251 X2.n1250 0.000932432
R4313 X2.n420 X2.n291 0.000932432
R4314 X2.n503 X2.n312 0.000932432
R4315 X2.n388 X2.n374 0.000898034
R4316 X2.n1079 X2.n1063 0.000898034
R4317 X2.n830 X2.n273 0.000875921
R4318 X2.n1127 X2.n151 0.000853808
R4319 X2.n745 X2.n529 0.000831695
R4320 X2.n533 X2.n532 0.000814286
R4321 X2.n912 X2.n911 0.000809582
R4322 X2.n996 X2.n200 0.000809582
R4323 X2.n681 X2.n680 0.000787469
R4324 X2.n650 X2.n649 0.000787469
R4325 X2.n424 X2.n423 0.000787469
R4326 X2.n512 X2.n511 0.000787469
R4327 X2.n1143 X2.n141 0.000765356
R4328 X2.n1201 X2.n116 0.000765356
R4329 X2.n1239 X2.n1238 0.000765356
R4330 X2.n1298 X2.n1297 0.000765356
R4331 X2.n742 X2.n531 0.000765356
R4332 X2.n1043 X2.n1042 0.000743243
R4333 X2.n863 X2.n259 0.00072113
R4334 X2.n716 X2.n20 0.000716216
R4335 X2.n613 X2.n49 0.000716216
R4336 X2.n829 X2.n270 0.000716216
R4337 X2.n1066 X2.n1065 0.000716216
R4338 X2.n874 X2.n873 0.000676904
R4339 X2.n549 X2.n548 0.000654791
R4340 X2.n611 X2.n598 0.000654791
R4341 X2.n1031 X2.n1030 0.000654791
R4342 X2.n1011 X2.n189 0.000588452
R4343 X2.n900 X2.n244 0.000566339
R4344 X2.n727 X2.n546 0.000522113
R4345 X2.n844 X2.n843 0.000522113
R4346 CLK_OUT.n1373 CLK_OUT 9.25617
R4347 CLK_OUT.n1374 CLK_OUT.n1373 9.23722
R4348 CLK_OUT.n1374 CLK_OUT 2.31448
R4349 CLK_OUT.n1344 CLK_OUT.n25 2.2505
R4350 CLK_OUT.n1346 CLK_OUT.n23 2.2505
R4351 CLK_OUT.n1350 CLK_OUT.n20 2.2505
R4352 CLK_OUT.n1352 CLK_OUT.n18 2.2505
R4353 CLK_OUT.n1356 CLK_OUT.n15 2.2505
R4354 CLK_OUT.n1358 CLK_OUT.n13 2.2505
R4355 CLK_OUT.n1362 CLK_OUT.n10 2.2505
R4356 CLK_OUT.n1363 CLK_OUT.n9 2.2505
R4357 CLK_OUT.n51 CLK_OUT.n6 2.2505
R4358 CLK_OUT.n1369 CLK_OUT.n4 2.2505
R4359 CLK_OUT.n1231 CLK_OUT.n2 2.2505
R4360 CLK_OUT.n64 CLK_OUT.n60 2.2505
R4361 CLK_OUT.n1206 CLK_OUT.n62 2.2505
R4362 CLK_OUT.n82 CLK_OUT.n72 2.2505
R4363 CLK_OUT.n1187 CLK_OUT.n74 2.2505
R4364 CLK_OUT.n957 CLK_OUT.n198 2.2505
R4365 CLK_OUT.n955 CLK_OUT.n200 2.2505
R4366 CLK_OUT.n951 CLK_OUT.n203 2.2505
R4367 CLK_OUT.n949 CLK_OUT.n205 2.2505
R4368 CLK_OUT.n945 CLK_OUT.n208 2.2505
R4369 CLK_OUT.n943 CLK_OUT.n210 2.2505
R4370 CLK_OUT.n939 CLK_OUT.n213 2.2505
R4371 CLK_OUT.n937 CLK_OUT.n215 2.2505
R4372 CLK_OUT.n361 CLK_OUT.n216 2.2505
R4373 CLK_OUT.n932 CLK_OUT.n219 2.2505
R4374 CLK_OUT.n617 CLK_OUT.n221 2.2505
R4375 CLK_OUT.n926 CLK_OUT.n224 2.2505
R4376 CLK_OUT.n664 CLK_OUT.n226 2.2505
R4377 CLK_OUT.n920 CLK_OUT.n229 2.2505
R4378 CLK_OUT.n320 CLK_OUT.n231 2.2505
R4379 CLK_OUT.n958 CLK_OUT.n957 2.2505
R4380 CLK_OUT.n955 CLK_OUT.n954 2.2505
R4381 CLK_OUT.n952 CLK_OUT.n951 2.2505
R4382 CLK_OUT.n949 CLK_OUT.n948 2.2505
R4383 CLK_OUT.n946 CLK_OUT.n945 2.2505
R4384 CLK_OUT.n943 CLK_OUT.n942 2.2505
R4385 CLK_OUT.n940 CLK_OUT.n939 2.2505
R4386 CLK_OUT.n937 CLK_OUT.n936 2.2505
R4387 CLK_OUT.n935 CLK_OUT.n216 2.2505
R4388 CLK_OUT.n932 CLK_OUT.n217 2.2505
R4389 CLK_OUT.n929 CLK_OUT.n221 2.2505
R4390 CLK_OUT.n926 CLK_OUT.n222 2.2505
R4391 CLK_OUT.n923 CLK_OUT.n226 2.2505
R4392 CLK_OUT.n920 CLK_OUT.n227 2.2505
R4393 CLK_OUT.n917 CLK_OUT.n231 2.2505
R4394 CLK_OUT.n1174 CLK_OUT.n1173 2.2505
R4395 CLK_OUT.n1175 CLK_OUT.n1171 2.2505
R4396 CLK_OUT.n1170 CLK_OUT.n95 2.2505
R4397 CLK_OUT.n1169 CLK_OUT.n1168 2.2505
R4398 CLK_OUT.n97 CLK_OUT.n96 2.2505
R4399 CLK_OUT.n1127 CLK_OUT.n1126 2.2505
R4400 CLK_OUT.n1134 CLK_OUT.n1125 2.2505
R4401 CLK_OUT.n1135 CLK_OUT.n1124 2.2505
R4402 CLK_OUT.n1123 CLK_OUT.n117 2.2505
R4403 CLK_OUT.n1122 CLK_OUT.n1121 2.2505
R4404 CLK_OUT.n119 CLK_OUT.n118 2.2505
R4405 CLK_OUT.n1100 CLK_OUT.n1099 2.2505
R4406 CLK_OUT.n1098 CLK_OUT.n130 2.2505
R4407 CLK_OUT.n1097 CLK_OUT.n1096 2.2505
R4408 CLK_OUT.n132 CLK_OUT.n131 2.2505
R4409 CLK_OUT.n1073 CLK_OUT.n1072 2.2505
R4410 CLK_OUT.n1074 CLK_OUT.n1071 2.2505
R4411 CLK_OUT.n1070 CLK_OUT.n143 2.2505
R4412 CLK_OUT.n1069 CLK_OUT.n1068 2.2505
R4413 CLK_OUT.n145 CLK_OUT.n144 2.2505
R4414 CLK_OUT.n1018 CLK_OUT.n1017 2.2505
R4415 CLK_OUT.n1019 CLK_OUT.n1016 2.2505
R4416 CLK_OUT.n1020 CLK_OUT.n1015 2.2505
R4417 CLK_OUT.n1021 CLK_OUT.n1014 2.2505
R4418 CLK_OUT.n1022 CLK_OUT.n1013 2.2505
R4419 CLK_OUT.n1012 CLK_OUT.n170 2.2505
R4420 CLK_OUT.n1011 CLK_OUT.n1010 2.2505
R4421 CLK_OUT.n172 CLK_OUT.n171 2.2505
R4422 CLK_OUT.n989 CLK_OUT.n988 2.2505
R4423 CLK_OUT.n987 CLK_OUT.n183 2.2505
R4424 CLK_OUT.n986 CLK_OUT.n985 2.2505
R4425 CLK_OUT.n185 CLK_OUT.n184 2.2505
R4426 CLK_OUT.n962 CLK_OUT.n961 2.2505
R4427 CLK_OUT.n963 CLK_OUT.n960 2.2505
R4428 CLK_OUT.n964 CLK_OUT.n963 2.2505
R4429 CLK_OUT.n962 CLK_OUT.n189 2.2505
R4430 CLK_OUT.n976 CLK_OUT.n185 2.2505
R4431 CLK_OUT.n985 CLK_OUT.n984 2.2505
R4432 CLK_OUT.n187 CLK_OUT.n183 2.2505
R4433 CLK_OUT.n990 CLK_OUT.n989 2.2505
R4434 CLK_OUT.n1001 CLK_OUT.n172 2.2505
R4435 CLK_OUT.n1010 CLK_OUT.n1009 2.2505
R4436 CLK_OUT.n170 CLK_OUT.n166 2.2505
R4437 CLK_OUT.n1023 CLK_OUT.n1022 2.2505
R4438 CLK_OUT.n1021 CLK_OUT.n159 2.2505
R4439 CLK_OUT.n1020 CLK_OUT.n157 2.2505
R4440 CLK_OUT.n1019 CLK_OUT.n155 2.2505
R4441 CLK_OUT.n1018 CLK_OUT.n153 2.2505
R4442 CLK_OUT.n1049 CLK_OUT.n145 2.2505
R4443 CLK_OUT.n1068 CLK_OUT.n1067 2.2505
R4444 CLK_OUT.n1060 CLK_OUT.n143 2.2505
R4445 CLK_OUT.n1075 CLK_OUT.n1074 2.2505
R4446 CLK_OUT.n1073 CLK_OUT.n136 2.2505
R4447 CLK_OUT.n1087 CLK_OUT.n132 2.2505
R4448 CLK_OUT.n1096 CLK_OUT.n1095 2.2505
R4449 CLK_OUT.n134 CLK_OUT.n130 2.2505
R4450 CLK_OUT.n1101 CLK_OUT.n1100 2.2505
R4451 CLK_OUT.n1112 CLK_OUT.n119 2.2505
R4452 CLK_OUT.n1121 CLK_OUT.n1120 2.2505
R4453 CLK_OUT.n117 CLK_OUT.n114 2.2505
R4454 CLK_OUT.n1136 CLK_OUT.n1135 2.2505
R4455 CLK_OUT.n1134 CLK_OUT.n1133 2.2505
R4456 CLK_OUT.n1127 CLK_OUT.n105 2.2505
R4457 CLK_OUT.n1149 CLK_OUT.n97 2.2505
R4458 CLK_OUT.n1168 CLK_OUT.n1167 2.2505
R4459 CLK_OUT.n1157 CLK_OUT.n95 2.2505
R4460 CLK_OUT.n1176 CLK_OUT.n1175 2.2505
R4461 CLK_OUT.n1174 CLK_OUT.n87 2.2505
R4462 CLK_OUT.n914 CLK_OUT.n234 2.2505
R4463 CLK_OUT.n913 CLK_OUT.n235 2.2505
R4464 CLK_OUT.n912 CLK_OUT.n236 2.2505
R4465 CLK_OUT.n733 CLK_OUT.n237 2.2505
R4466 CLK_OUT.n908 CLK_OUT.n239 2.2505
R4467 CLK_OUT.n907 CLK_OUT.n240 2.2505
R4468 CLK_OUT.n906 CLK_OUT.n241 2.2505
R4469 CLK_OUT.n748 CLK_OUT.n242 2.2505
R4470 CLK_OUT.n902 CLK_OUT.n244 2.2505
R4471 CLK_OUT.n901 CLK_OUT.n245 2.2505
R4472 CLK_OUT.n900 CLK_OUT.n246 2.2505
R4473 CLK_OUT.n298 CLK_OUT.n247 2.2505
R4474 CLK_OUT.n896 CLK_OUT.n249 2.2505
R4475 CLK_OUT.n895 CLK_OUT.n250 2.2505
R4476 CLK_OUT.n894 CLK_OUT.n251 2.2505
R4477 CLK_OUT.n787 CLK_OUT.n252 2.2505
R4478 CLK_OUT.n890 CLK_OUT.n254 2.2505
R4479 CLK_OUT.n889 CLK_OUT.n255 2.2505
R4480 CLK_OUT.n888 CLK_OUT.n256 2.2505
R4481 CLK_OUT.n805 CLK_OUT.n257 2.2505
R4482 CLK_OUT.n884 CLK_OUT.n259 2.2505
R4483 CLK_OUT.n883 CLK_OUT.n260 2.2505
R4484 CLK_OUT.n882 CLK_OUT.n261 2.2505
R4485 CLK_OUT.n822 CLK_OUT.n262 2.2505
R4486 CLK_OUT.n878 CLK_OUT.n264 2.2505
R4487 CLK_OUT.n877 CLK_OUT.n265 2.2505
R4488 CLK_OUT.n876 CLK_OUT.n266 2.2505
R4489 CLK_OUT.n281 CLK_OUT.n267 2.2505
R4490 CLK_OUT.n872 CLK_OUT.n269 2.2505
R4491 CLK_OUT.n871 CLK_OUT.n270 2.2505
R4492 CLK_OUT.n870 CLK_OUT.n271 2.2505
R4493 CLK_OUT.n867 CLK_OUT.n866 2.2505
R4494 CLK_OUT.n275 CLK_OUT.n28 2.2505
R4495 CLK_OUT.n1340 CLK_OUT.n1339 2.2505
R4496 CLK_OUT.n1341 CLK_OUT.n1340 2.2505
R4497 CLK_OUT.n28 CLK_OUT.n27 2.2505
R4498 CLK_OUT.n868 CLK_OUT.n867 2.2505
R4499 CLK_OUT.n870 CLK_OUT.n869 2.2505
R4500 CLK_OUT.n871 CLK_OUT.n268 2.2505
R4501 CLK_OUT.n873 CLK_OUT.n872 2.2505
R4502 CLK_OUT.n874 CLK_OUT.n267 2.2505
R4503 CLK_OUT.n876 CLK_OUT.n875 2.2505
R4504 CLK_OUT.n877 CLK_OUT.n263 2.2505
R4505 CLK_OUT.n879 CLK_OUT.n878 2.2505
R4506 CLK_OUT.n880 CLK_OUT.n262 2.2505
R4507 CLK_OUT.n882 CLK_OUT.n881 2.2505
R4508 CLK_OUT.n883 CLK_OUT.n258 2.2505
R4509 CLK_OUT.n885 CLK_OUT.n884 2.2505
R4510 CLK_OUT.n886 CLK_OUT.n257 2.2505
R4511 CLK_OUT.n888 CLK_OUT.n887 2.2505
R4512 CLK_OUT.n889 CLK_OUT.n253 2.2505
R4513 CLK_OUT.n891 CLK_OUT.n890 2.2505
R4514 CLK_OUT.n892 CLK_OUT.n252 2.2505
R4515 CLK_OUT.n894 CLK_OUT.n893 2.2505
R4516 CLK_OUT.n895 CLK_OUT.n248 2.2505
R4517 CLK_OUT.n897 CLK_OUT.n896 2.2505
R4518 CLK_OUT.n898 CLK_OUT.n247 2.2505
R4519 CLK_OUT.n900 CLK_OUT.n899 2.2505
R4520 CLK_OUT.n901 CLK_OUT.n243 2.2505
R4521 CLK_OUT.n903 CLK_OUT.n902 2.2505
R4522 CLK_OUT.n904 CLK_OUT.n242 2.2505
R4523 CLK_OUT.n906 CLK_OUT.n905 2.2505
R4524 CLK_OUT.n907 CLK_OUT.n238 2.2505
R4525 CLK_OUT.n909 CLK_OUT.n908 2.2505
R4526 CLK_OUT.n910 CLK_OUT.n237 2.2505
R4527 CLK_OUT.n912 CLK_OUT.n911 2.2505
R4528 CLK_OUT.n913 CLK_OUT.n233 2.2505
R4529 CLK_OUT.n915 CLK_OUT.n914 2.2505
R4530 CLK_OUT.n1344 CLK_OUT.n1343 2.2505
R4531 CLK_OUT.n1347 CLK_OUT.n1346 2.2505
R4532 CLK_OUT.n1350 CLK_OUT.n1349 2.2505
R4533 CLK_OUT.n1353 CLK_OUT.n1352 2.2505
R4534 CLK_OUT.n1356 CLK_OUT.n1355 2.2505
R4535 CLK_OUT.n1359 CLK_OUT.n1358 2.2505
R4536 CLK_OUT.n1362 CLK_OUT.n1361 2.2505
R4537 CLK_OUT.n1363 CLK_OUT.n7 2.2505
R4538 CLK_OUT.n1366 CLK_OUT.n6 2.2505
R4539 CLK_OUT.n1369 CLK_OUT.n1 2.2505
R4540 CLK_OUT.n1220 CLK_OUT.n60 2.2505
R4541 CLK_OUT.n62 CLK_OUT.n61 2.2505
R4542 CLK_OUT.n1200 CLK_OUT.n72 2.2505
R4543 CLK_OUT.n74 CLK_OUT.n73 2.2505
R4544 CLK_OUT.n2 CLK_OUT.n0 2.2505
R4545 CLK_OUT.n31 CLK_OUT.n30 2.2005
R4546 CLK_OUT.n1186 CLK_OUT.n86 2.2005
R4547 CLK_OUT.n1189 CLK_OUT.n1188 2.2005
R4548 CLK_OUT.n77 CLK_OUT.n75 2.2005
R4549 CLK_OUT.n1196 CLK_OUT.n1195 2.2005
R4550 CLK_OUT.n1194 CLK_OUT.n76 2.2005
R4551 CLK_OUT.n84 CLK_OUT.n83 2.2005
R4552 CLK_OUT.n81 CLK_OUT.n80 2.2005
R4553 CLK_OUT.n78 CLK_OUT.n71 2.2005
R4554 CLK_OUT.n1204 CLK_OUT.n68 2.2005
R4555 CLK_OUT.n1208 CLK_OUT.n1207 2.2005
R4556 CLK_OUT.n1205 CLK_OUT.n70 2.2005
R4557 CLK_OUT.n69 CLK_OUT.n63 2.2005
R4558 CLK_OUT.n1216 CLK_OUT.n1215 2.2005
R4559 CLK_OUT.n1214 CLK_OUT.n65 2.2005
R4560 CLK_OUT.n59 CLK_OUT.n58 2.2005
R4561 CLK_OUT.n1225 CLK_OUT.n1224 2.2005
R4562 CLK_OUT.n1227 CLK_OUT.n57 2.2005
R4563 CLK_OUT.n1229 CLK_OUT.n1228 2.2005
R4564 CLK_OUT.n1230 CLK_OUT.n56 2.2005
R4565 CLK_OUT.n1234 CLK_OUT.n1233 2.2005
R4566 CLK_OUT.n1232 CLK_OUT.n54 2.2005
R4567 CLK_OUT.n1240 CLK_OUT.n1239 2.2005
R4568 CLK_OUT.n1242 CLK_OUT.n1241 2.2005
R4569 CLK_OUT.n1245 CLK_OUT.n1244 2.2005
R4570 CLK_OUT.n1247 CLK_OUT.n1246 2.2005
R4571 CLK_OUT.n1250 CLK_OUT.n1249 2.2005
R4572 CLK_OUT.n1248 CLK_OUT.n52 2.2005
R4573 CLK_OUT.n1256 CLK_OUT.n1255 2.2005
R4574 CLK_OUT.n1257 CLK_OUT.n50 2.2005
R4575 CLK_OUT.n1259 CLK_OUT.n1258 2.2005
R4576 CLK_OUT.n1261 CLK_OUT.n1260 2.2005
R4577 CLK_OUT.n1263 CLK_OUT.n1262 2.2005
R4578 CLK_OUT.n1265 CLK_OUT.n1264 2.2005
R4579 CLK_OUT.n1267 CLK_OUT.n1266 2.2005
R4580 CLK_OUT.n48 CLK_OUT.n47 2.2005
R4581 CLK_OUT.n1273 CLK_OUT.n1272 2.2005
R4582 CLK_OUT.n1275 CLK_OUT.n46 2.2005
R4583 CLK_OUT.n1277 CLK_OUT.n1276 2.2005
R4584 CLK_OUT.n1280 CLK_OUT.n1279 2.2005
R4585 CLK_OUT.n1282 CLK_OUT.n1281 2.2005
R4586 CLK_OUT.n1285 CLK_OUT.n1284 2.2005
R4587 CLK_OUT.n1283 CLK_OUT.n44 2.2005
R4588 CLK_OUT.n1291 CLK_OUT.n1290 2.2005
R4589 CLK_OUT.n1292 CLK_OUT.n43 2.2005
R4590 CLK_OUT.n1295 CLK_OUT.n1294 2.2005
R4591 CLK_OUT.n1297 CLK_OUT.n42 2.2005
R4592 CLK_OUT.n1299 CLK_OUT.n1298 2.2005
R4593 CLK_OUT.n1302 CLK_OUT.n1301 2.2005
R4594 CLK_OUT.n1300 CLK_OUT.n40 2.2005
R4595 CLK_OUT.n1310 CLK_OUT.n1309 2.2005
R4596 CLK_OUT.n1312 CLK_OUT.n1311 2.2005
R4597 CLK_OUT.n1314 CLK_OUT.n1313 2.2005
R4598 CLK_OUT.n1316 CLK_OUT.n1315 2.2005
R4599 CLK_OUT.n1318 CLK_OUT.n1317 2.2005
R4600 CLK_OUT.n1320 CLK_OUT.n1319 2.2005
R4601 CLK_OUT.n1323 CLK_OUT.n1322 2.2005
R4602 CLK_OUT.n1324 CLK_OUT.n36 2.2005
R4603 CLK_OUT.n1326 CLK_OUT.n1325 2.2005
R4604 CLK_OUT.n1328 CLK_OUT.n1327 2.2005
R4605 CLK_OUT.n1330 CLK_OUT.n1329 2.2005
R4606 CLK_OUT.n712 CLK_OUT.n711 2.2005
R4607 CLK_OUT.n700 CLK_OUT.n699 2.2005
R4608 CLK_OUT.n698 CLK_OUT.n697 2.2005
R4609 CLK_OUT.n691 CLK_OUT.n690 2.2005
R4610 CLK_OUT.n689 CLK_OUT.n688 2.2005
R4611 CLK_OUT.n682 CLK_OUT.n327 2.2005
R4612 CLK_OUT.n673 CLK_OUT.n331 2.2005
R4613 CLK_OUT.n675 CLK_OUT.n674 2.2005
R4614 CLK_OUT.n665 CLK_OUT.n333 2.2005
R4615 CLK_OUT.n667 CLK_OUT.n666 2.2005
R4616 CLK_OUT.n663 CLK_OUT.n662 2.2005
R4617 CLK_OUT.n655 CLK_OUT.n336 2.2005
R4618 CLK_OUT.n649 CLK_OUT.n648 2.2005
R4619 CLK_OUT.n647 CLK_OUT.n646 2.2005
R4620 CLK_OUT.n642 CLK_OUT.n641 2.2005
R4621 CLK_OUT.n640 CLK_OUT.n639 2.2005
R4622 CLK_OUT.n634 CLK_OUT.n633 2.2005
R4623 CLK_OUT.n632 CLK_OUT.n631 2.2005
R4624 CLK_OUT.n625 CLK_OUT.n348 2.2005
R4625 CLK_OUT.n619 CLK_OUT.n618 2.2005
R4626 CLK_OUT.n616 CLK_OUT.n615 2.2005
R4627 CLK_OUT.n606 CLK_OUT.n353 2.2005
R4628 CLK_OUT.n608 CLK_OUT.n607 2.2005
R4629 CLK_OUT.n601 CLK_OUT.n600 2.2005
R4630 CLK_OUT.n599 CLK_OUT.n598 2.2005
R4631 CLK_OUT.n592 CLK_OUT.n591 2.2005
R4632 CLK_OUT.n590 CLK_OUT.n589 2.2005
R4633 CLK_OUT.n583 CLK_OUT.n582 2.2005
R4634 CLK_OUT.n581 CLK_OUT.n580 2.2005
R4635 CLK_OUT.n574 CLK_OUT.n573 2.2005
R4636 CLK_OUT.n572 CLK_OUT.n571 2.2005
R4637 CLK_OUT.n565 CLK_OUT.n564 2.2005
R4638 CLK_OUT.n563 CLK_OUT.n562 2.2005
R4639 CLK_OUT.n557 CLK_OUT.n372 2.2005
R4640 CLK_OUT.n548 CLK_OUT.n376 2.2005
R4641 CLK_OUT.n550 CLK_OUT.n549 2.2005
R4642 CLK_OUT.n546 CLK_OUT.n545 2.2005
R4643 CLK_OUT.n538 CLK_OUT.n379 2.2005
R4644 CLK_OUT.n532 CLK_OUT.n531 2.2005
R4645 CLK_OUT.n530 CLK_OUT.n529 2.2005
R4646 CLK_OUT.n525 CLK_OUT.n524 2.2005
R4647 CLK_OUT.n523 CLK_OUT.n522 2.2005
R4648 CLK_OUT.n517 CLK_OUT.n516 2.2005
R4649 CLK_OUT.n515 CLK_OUT.n514 2.2005
R4650 CLK_OUT.n508 CLK_OUT.n391 2.2005
R4651 CLK_OUT.n502 CLK_OUT.n501 2.2005
R4652 CLK_OUT.n499 CLK_OUT.n498 2.2005
R4653 CLK_OUT.n489 CLK_OUT.n396 2.2005
R4654 CLK_OUT.n491 CLK_OUT.n490 2.2005
R4655 CLK_OUT.n484 CLK_OUT.n483 2.2005
R4656 CLK_OUT.n482 CLK_OUT.n481 2.2005
R4657 CLK_OUT.n475 CLK_OUT.n474 2.2005
R4658 CLK_OUT.n473 CLK_OUT.n472 2.2005
R4659 CLK_OUT.n466 CLK_OUT.n465 2.2005
R4660 CLK_OUT.n464 CLK_OUT.n463 2.2005
R4661 CLK_OUT.n458 CLK_OUT.n457 2.2005
R4662 CLK_OUT.n456 CLK_OUT.n455 2.2005
R4663 CLK_OUT.n449 CLK_OUT.n411 2.2005
R4664 CLK_OUT.n440 CLK_OUT.n415 2.2005
R4665 CLK_OUT.n442 CLK_OUT.n441 2.2005
R4666 CLK_OUT.n435 CLK_OUT.n434 2.2005
R4667 CLK_OUT.n421 CLK_OUT.n195 2.2005
R4668 CLK_OUT.n965 CLK_OUT.n194 2.2005
R4669 CLK_OUT.n967 CLK_OUT.n966 2.2005
R4670 CLK_OUT.n974 CLK_OUT.n973 2.2005
R4671 CLK_OUT.n975 CLK_OUT.n188 2.2005
R4672 CLK_OUT.n978 CLK_OUT.n977 2.2005
R4673 CLK_OUT.n980 CLK_OUT.n186 2.2005
R4674 CLK_OUT.n983 CLK_OUT.n982 2.2005
R4675 CLK_OUT.n182 CLK_OUT.n181 2.2005
R4676 CLK_OUT.n993 CLK_OUT.n991 2.2005
R4677 CLK_OUT.n177 CLK_OUT.n176 2.2005
R4678 CLK_OUT.n1000 CLK_OUT.n999 2.2005
R4679 CLK_OUT.n1003 CLK_OUT.n1002 2.2005
R4680 CLK_OUT.n1005 CLK_OUT.n173 2.2005
R4681 CLK_OUT.n1008 CLK_OUT.n1007 2.2005
R4682 CLK_OUT.n174 CLK_OUT.n164 2.2005
R4683 CLK_OUT.n1026 CLK_OUT.n1025 2.2005
R4684 CLK_OUT.n1024 CLK_OUT.n165 2.2005
R4685 CLK_OUT.n169 CLK_OUT.n168 2.2005
R4686 CLK_OUT.n167 CLK_OUT.n160 2.2005
R4687 CLK_OUT.n1034 CLK_OUT.n1033 2.2005
R4688 CLK_OUT.n1036 CLK_OUT.n1035 2.2005
R4689 CLK_OUT.n1038 CLK_OUT.n1037 2.2005
R4690 CLK_OUT.n1040 CLK_OUT.n1039 2.2005
R4691 CLK_OUT.n1042 CLK_OUT.n1041 2.2005
R4692 CLK_OUT.n1044 CLK_OUT.n1043 2.2005
R4693 CLK_OUT.n1047 CLK_OUT.n1046 2.2005
R4694 CLK_OUT.n1048 CLK_OUT.n152 2.2005
R4695 CLK_OUT.n1052 CLK_OUT.n1050 2.2005
R4696 CLK_OUT.n148 CLK_OUT.n146 2.2005
R4697 CLK_OUT.n1066 CLK_OUT.n1065 2.2005
R4698 CLK_OUT.n1064 CLK_OUT.n147 2.2005
R4699 CLK_OUT.n1062 CLK_OUT.n1061 2.2005
R4700 CLK_OUT.n1058 CLK_OUT.n142 2.2005
R4701 CLK_OUT.n1076 CLK_OUT.n141 2.2005
R4702 CLK_OUT.n1078 CLK_OUT.n1077 2.2005
R4703 CLK_OUT.n1085 CLK_OUT.n1084 2.2005
R4704 CLK_OUT.n1086 CLK_OUT.n135 2.2005
R4705 CLK_OUT.n1089 CLK_OUT.n1088 2.2005
R4706 CLK_OUT.n1091 CLK_OUT.n133 2.2005
R4707 CLK_OUT.n1094 CLK_OUT.n1093 2.2005
R4708 CLK_OUT.n129 CLK_OUT.n128 2.2005
R4709 CLK_OUT.n1104 CLK_OUT.n1102 2.2005
R4710 CLK_OUT.n124 CLK_OUT.n123 2.2005
R4711 CLK_OUT.n1111 CLK_OUT.n1110 2.2005
R4712 CLK_OUT.n1114 CLK_OUT.n1113 2.2005
R4713 CLK_OUT.n1116 CLK_OUT.n120 2.2005
R4714 CLK_OUT.n1119 CLK_OUT.n1118 2.2005
R4715 CLK_OUT.n121 CLK_OUT.n112 2.2005
R4716 CLK_OUT.n1139 CLK_OUT.n1138 2.2005
R4717 CLK_OUT.n1137 CLK_OUT.n113 2.2005
R4718 CLK_OUT.n116 CLK_OUT.n115 2.2005
R4719 CLK_OUT.n1129 CLK_OUT.n1128 2.2005
R4720 CLK_OUT.n1132 CLK_OUT.n1131 2.2005
R4721 CLK_OUT.n1130 CLK_OUT.n106 2.2005
R4722 CLK_OUT.n1147 CLK_OUT.n1146 2.2005
R4723 CLK_OUT.n1148 CLK_OUT.n104 2.2005
R4724 CLK_OUT.n1151 CLK_OUT.n1150 2.2005
R4725 CLK_OUT.n102 CLK_OUT.n98 2.2005
R4726 CLK_OUT.n1166 CLK_OUT.n1165 2.2005
R4727 CLK_OUT.n101 CLK_OUT.n99 2.2005
R4728 CLK_OUT.n1159 CLK_OUT.n1158 2.2005
R4729 CLK_OUT.n94 CLK_OUT.n92 2.2005
R4730 CLK_OUT.n1179 CLK_OUT.n1178 2.2005
R4731 CLK_OUT.n1177 CLK_OUT.n93 2.2005
R4732 CLK_OUT.n714 CLK_OUT.n713 2.2005
R4733 CLK_OUT.n723 CLK_OUT.n722 2.2005
R4734 CLK_OUT.n725 CLK_OUT.n724 2.2005
R4735 CLK_OUT.n727 CLK_OUT.n726 2.2005
R4736 CLK_OUT.n729 CLK_OUT.n728 2.2005
R4737 CLK_OUT.n730 CLK_OUT.n307 2.2005
R4738 CLK_OUT.n732 CLK_OUT.n731 2.2005
R4739 CLK_OUT.n735 CLK_OUT.n734 2.2005
R4740 CLK_OUT.n737 CLK_OUT.n736 2.2005
R4741 CLK_OUT.n739 CLK_OUT.n738 2.2005
R4742 CLK_OUT.n741 CLK_OUT.n740 2.2005
R4743 CLK_OUT.n743 CLK_OUT.n742 2.2005
R4744 CLK_OUT.n744 CLK_OUT.n303 2.2005
R4745 CLK_OUT.n747 CLK_OUT.n746 2.2005
R4746 CLK_OUT.n749 CLK_OUT.n302 2.2005
R4747 CLK_OUT.n751 CLK_OUT.n750 2.2005
R4748 CLK_OUT.n754 CLK_OUT.n753 2.2005
R4749 CLK_OUT.n752 CLK_OUT.n300 2.2005
R4750 CLK_OUT.n762 CLK_OUT.n761 2.2005
R4751 CLK_OUT.n764 CLK_OUT.n763 2.2005
R4752 CLK_OUT.n766 CLK_OUT.n765 2.2005
R4753 CLK_OUT.n768 CLK_OUT.n767 2.2005
R4754 CLK_OUT.n770 CLK_OUT.n769 2.2005
R4755 CLK_OUT.n772 CLK_OUT.n771 2.2005
R4756 CLK_OUT.n774 CLK_OUT.n773 2.2005
R4757 CLK_OUT.n776 CLK_OUT.n775 2.2005
R4758 CLK_OUT.n778 CLK_OUT.n777 2.2005
R4759 CLK_OUT.n780 CLK_OUT.n779 2.2005
R4760 CLK_OUT.n294 CLK_OUT.n293 2.2005
R4761 CLK_OUT.n786 CLK_OUT.n785 2.2005
R4762 CLK_OUT.n788 CLK_OUT.n292 2.2005
R4763 CLK_OUT.n790 CLK_OUT.n789 2.2005
R4764 CLK_OUT.n792 CLK_OUT.n791 2.2005
R4765 CLK_OUT.n794 CLK_OUT.n793 2.2005
R4766 CLK_OUT.n796 CLK_OUT.n795 2.2005
R4767 CLK_OUT.n798 CLK_OUT.n797 2.2005
R4768 CLK_OUT.n290 CLK_OUT.n289 2.2005
R4769 CLK_OUT.n804 CLK_OUT.n803 2.2005
R4770 CLK_OUT.n806 CLK_OUT.n288 2.2005
R4771 CLK_OUT.n808 CLK_OUT.n807 2.2005
R4772 CLK_OUT.n811 CLK_OUT.n810 2.2005
R4773 CLK_OUT.n813 CLK_OUT.n812 2.2005
R4774 CLK_OUT.n815 CLK_OUT.n814 2.2005
R4775 CLK_OUT.n286 CLK_OUT.n285 2.2005
R4776 CLK_OUT.n821 CLK_OUT.n820 2.2005
R4777 CLK_OUT.n823 CLK_OUT.n284 2.2005
R4778 CLK_OUT.n825 CLK_OUT.n824 2.2005
R4779 CLK_OUT.n828 CLK_OUT.n827 2.2005
R4780 CLK_OUT.n830 CLK_OUT.n829 2.2005
R4781 CLK_OUT.n833 CLK_OUT.n832 2.2005
R4782 CLK_OUT.n831 CLK_OUT.n282 2.2005
R4783 CLK_OUT.n840 CLK_OUT.n839 2.2005
R4784 CLK_OUT.n842 CLK_OUT.n841 2.2005
R4785 CLK_OUT.n844 CLK_OUT.n843 2.2005
R4786 CLK_OUT.n846 CLK_OUT.n845 2.2005
R4787 CLK_OUT.n848 CLK_OUT.n847 2.2005
R4788 CLK_OUT.n850 CLK_OUT.n849 2.2005
R4789 CLK_OUT.n855 CLK_OUT.n851 2.2005
R4790 CLK_OUT.n857 CLK_OUT.n856 2.2005
R4791 CLK_OUT.n854 CLK_OUT.n853 2.2005
R4792 CLK_OUT.n852 CLK_OUT.n272 2.2005
R4793 CLK_OUT.n865 CLK_OUT.n864 2.2005
R4794 CLK_OUT.n863 CLK_OUT.n273 2.2005
R4795 CLK_OUT.n277 CLK_OUT.n276 2.2005
R4796 CLK_OUT.n32 CLK_OUT.n29 2.2005
R4797 CLK_OUT.n1345 CLK_OUT.n24 1.8005
R4798 CLK_OUT.n38 CLK_OUT.n21 1.8005
R4799 CLK_OUT.n1351 CLK_OUT.n19 1.8005
R4800 CLK_OUT.n1296 CLK_OUT.n16 1.8005
R4801 CLK_OUT.n1357 CLK_OUT.n14 1.8005
R4802 CLK_OUT.n1274 CLK_OUT.n11 1.8005
R4803 CLK_OUT.n1364 CLK_OUT.n8 1.8005
R4804 CLK_OUT.n1368 CLK_OUT.n5 1.8005
R4805 CLK_OUT.n1370 CLK_OUT.n3 1.8005
R4806 CLK_OUT.n1223 CLK_OUT.n1222 1.8005
R4807 CLK_OUT.n1218 CLK_OUT.n1217 1.8005
R4808 CLK_OUT.n1203 CLK_OUT.n1202 1.8005
R4809 CLK_OUT.n1198 CLK_OUT.n1197 1.8005
R4810 CLK_OUT.n956 CLK_OUT.n199 1.8005
R4811 CLK_OUT.n404 CLK_OUT.n201 1.8005
R4812 CLK_OUT.n950 CLK_OUT.n204 1.8005
R4813 CLK_OUT.n500 CLK_OUT.n206 1.8005
R4814 CLK_OUT.n944 CLK_OUT.n209 1.8005
R4815 CLK_OUT.n547 CLK_OUT.n211 1.8005
R4816 CLK_OUT.n938 CLK_OUT.n214 1.8005
R4817 CLK_OUT.n933 CLK_OUT.n218 1.8005
R4818 CLK_OUT.n931 CLK_OUT.n220 1.8005
R4819 CLK_OUT.n927 CLK_OUT.n223 1.8005
R4820 CLK_OUT.n925 CLK_OUT.n225 1.8005
R4821 CLK_OUT.n921 CLK_OUT.n228 1.8005
R4822 CLK_OUT.n919 CLK_OUT.n230 1.8005
R4823 CLK_OUT.n956 CLK_OUT.n197 1.8005
R4824 CLK_OUT.n953 CLK_OUT.n201 1.8005
R4825 CLK_OUT.n950 CLK_OUT.n202 1.8005
R4826 CLK_OUT.n947 CLK_OUT.n206 1.8005
R4827 CLK_OUT.n944 CLK_OUT.n207 1.8005
R4828 CLK_OUT.n941 CLK_OUT.n211 1.8005
R4829 CLK_OUT.n938 CLK_OUT.n212 1.8005
R4830 CLK_OUT.n934 CLK_OUT.n933 1.8005
R4831 CLK_OUT.n931 CLK_OUT.n930 1.8005
R4832 CLK_OUT.n928 CLK_OUT.n927 1.8005
R4833 CLK_OUT.n925 CLK_OUT.n924 1.8005
R4834 CLK_OUT.n922 CLK_OUT.n921 1.8005
R4835 CLK_OUT.n919 CLK_OUT.n918 1.8005
R4836 CLK_OUT.n1172 CLK_OUT.n88 1.8005
R4837 CLK_OUT.n1185 CLK_OUT.n88 1.8005
R4838 CLK_OUT.n1338 CLK_OUT.n26 1.8005
R4839 CLK_OUT.n1342 CLK_OUT.n26 1.8005
R4840 CLK_OUT.n1345 CLK_OUT.n22 1.8005
R4841 CLK_OUT.n1348 CLK_OUT.n21 1.8005
R4842 CLK_OUT.n1351 CLK_OUT.n17 1.8005
R4843 CLK_OUT.n1354 CLK_OUT.n16 1.8005
R4844 CLK_OUT.n1357 CLK_OUT.n12 1.8005
R4845 CLK_OUT.n1360 CLK_OUT.n11 1.8005
R4846 CLK_OUT.n1365 CLK_OUT.n1364 1.8005
R4847 CLK_OUT.n1368 CLK_OUT.n1367 1.8005
R4848 CLK_OUT.n1371 CLK_OUT.n1370 1.8005
R4849 CLK_OUT.n1222 CLK_OUT.n1221 1.8005
R4850 CLK_OUT.n1219 CLK_OUT.n1218 1.8005
R4851 CLK_OUT.n1202 CLK_OUT.n1201 1.8005
R4852 CLK_OUT.n1199 CLK_OUT.n1198 1.8005
R4853 CLK_OUT.n959 CLK_OUT.n196 1.5005
R4854 CLK_OUT.n433 CLK_OUT.n196 1.5005
R4855 CLK_OUT.n715 CLK_OUT.n232 1.5005
R4856 CLK_OUT.n916 CLK_OUT.n232 1.5005
R4857 CLK_OUT.n719 CLK_OUT.n315 1.1125
R4858 CLK_OUT.n1164 CLK_OUT.n1163 1.10836
R4859 CLK_OUT.n1156 CLK_OUT.n100 1.10443
R4860 CLK_OUT.n1182 CLK_OUT.n90 1.10381
R4861 CLK_OUT.n718 CLK_OUT.n316 1.10372
R4862 CLK_OUT.n1152 CLK_OUT.n103 1.10339
R4863 CLK_OUT.n1159 CLK_OUT.n91 1.10272
R4864 CLK_OUT.n1162 CLK_OUT.n101 1.10272
R4865 CLK_OUT.n1155 CLK_OUT.n102 1.10272
R4866 CLK_OUT.n722 CLK_OUT.n721 1.10263
R4867 CLK_OUT.n725 CLK_OUT.n314 1.10263
R4868 CLK_OUT.n1332 CLK_OUT.n1331 1.1005
R4869 CLK_OUT.n1191 CLK_OUT.n1190 1.1005
R4870 CLK_OUT.n1193 CLK_OUT.n1192 1.1005
R4871 CLK_OUT.n79 CLK_OUT.n67 1.1005
R4872 CLK_OUT.n1210 CLK_OUT.n1209 1.1005
R4873 CLK_OUT.n1211 CLK_OUT.n66 1.1005
R4874 CLK_OUT.n1213 CLK_OUT.n1212 1.1005
R4875 CLK_OUT.n1226 CLK_OUT.n55 1.1005
R4876 CLK_OUT.n1236 CLK_OUT.n1235 1.1005
R4877 CLK_OUT.n1238 CLK_OUT.n1237 1.1005
R4878 CLK_OUT.n1243 CLK_OUT.n53 1.1005
R4879 CLK_OUT.n1252 CLK_OUT.n1251 1.1005
R4880 CLK_OUT.n1254 CLK_OUT.n1253 1.1005
R4881 CLK_OUT.n1260 CLK_OUT.n49 1.1005
R4882 CLK_OUT.n1269 CLK_OUT.n1268 1.1005
R4883 CLK_OUT.n1271 CLK_OUT.n1270 1.1005
R4884 CLK_OUT.n1278 CLK_OUT.n45 1.1005
R4885 CLK_OUT.n1287 CLK_OUT.n1286 1.1005
R4886 CLK_OUT.n1289 CLK_OUT.n1288 1.1005
R4887 CLK_OUT.n1293 CLK_OUT.n41 1.1005
R4888 CLK_OUT.n1304 CLK_OUT.n1303 1.1005
R4889 CLK_OUT.n1308 CLK_OUT.n1307 1.1005
R4890 CLK_OUT.n1306 CLK_OUT.n39 1.1005
R4891 CLK_OUT.n1305 CLK_OUT.n37 1.1005
R4892 CLK_OUT.n1321 CLK_OUT.n35 1.1005
R4893 CLK_OUT.n89 CLK_OUT.n85 1.1005
R4894 CLK_OUT.n968 CLK_OUT.n192 1.1005
R4895 CLK_OUT.n994 CLK_OUT.n179 1.1005
R4896 CLK_OUT.n1053 CLK_OUT.n150 1.1005
R4897 CLK_OUT.n1079 CLK_OUT.n139 1.1005
R4898 CLK_OUT.n1105 CLK_OUT.n126 1.1005
R4899 CLK_OUT.n1181 CLK_OUT.n1180 1.1005
R4900 CLK_OUT.n1161 CLK_OUT.n1160 1.1005
R4901 CLK_OUT.n1154 CLK_OUT.n1153 1.1005
R4902 CLK_OUT.n1145 CLK_OUT.n1144 1.1005
R4903 CLK_OUT.n1141 CLK_OUT.n1140 1.1005
R4904 CLK_OUT.n1107 CLK_OUT.n1106 1.1005
R4905 CLK_OUT.n1083 CLK_OUT.n1082 1.1005
R4906 CLK_OUT.n1081 CLK_OUT.n1080 1.1005
R4907 CLK_OUT.n1057 CLK_OUT.n1056 1.1005
R4908 CLK_OUT.n1055 CLK_OUT.n1054 1.1005
R4909 CLK_OUT.n1030 CLK_OUT.n156 1.1005
R4910 CLK_OUT.n1028 CLK_OUT.n1027 1.1005
R4911 CLK_OUT.n996 CLK_OUT.n995 1.1005
R4912 CLK_OUT.n972 CLK_OUT.n971 1.1005
R4913 CLK_OUT.n970 CLK_OUT.n969 1.1005
R4914 CLK_OUT.n430 CLK_OUT.n423 1.1005
R4915 CLK_OUT.n429 CLK_OUT.n420 1.1005
R4916 CLK_OUT.n422 CLK_OUT.n193 1.1005
R4917 CLK_OUT.n432 CLK_OUT.n431 1.1005
R4918 CLK_OUT.n711 CLK_OUT.n710 1.1005
R4919 CLK_OUT.n702 CLK_OUT.n701 1.1005
R4920 CLK_OUT.n700 CLK_OUT.n322 1.1005
R4921 CLK_OUT.n697 CLK_OUT.n696 1.1005
R4922 CLK_OUT.n693 CLK_OUT.n692 1.1005
R4923 CLK_OUT.n686 CLK_OUT.n329 1.1005
R4924 CLK_OUT.n688 CLK_OUT.n687 1.1005
R4925 CLK_OUT.n685 CLK_OUT.n328 1.1005
R4926 CLK_OUT.n680 CLK_OUT.n679 1.1005
R4927 CLK_OUT.n669 CLK_OUT.n668 1.1005
R4928 CLK_OUT.n667 CLK_OUT.n334 1.1005
R4929 CLK_OUT.n659 CLK_OUT.n335 1.1005
R4930 CLK_OUT.n657 CLK_OUT.n656 1.1005
R4931 CLK_OUT.n655 CLK_OUT.n338 1.1005
R4932 CLK_OUT.n654 CLK_OUT.n653 1.1005
R4933 CLK_OUT.n341 CLK_OUT.n340 1.1005
R4934 CLK_OUT.n636 CLK_OUT.n345 1.1005
R4935 CLK_OUT.n635 CLK_OUT.n634 1.1005
R4936 CLK_OUT.n347 CLK_OUT.n346 1.1005
R4937 CLK_OUT.n627 CLK_OUT.n626 1.1005
R4938 CLK_OUT.n625 CLK_OUT.n350 1.1005
R4939 CLK_OUT.n624 CLK_OUT.n623 1.1005
R4940 CLK_OUT.n621 CLK_OUT.n620 1.1005
R4941 CLK_OUT.n615 CLK_OUT.n352 1.1005
R4942 CLK_OUT.n612 CLK_OUT.n353 1.1005
R4943 CLK_OUT.n609 CLK_OUT.n354 1.1005
R4944 CLK_OUT.n603 CLK_OUT.n355 1.1005
R4945 CLK_OUT.n602 CLK_OUT.n601 1.1005
R4946 CLK_OUT.n357 CLK_OUT.n356 1.1005
R4947 CLK_OUT.n594 CLK_OUT.n593 1.1005
R4948 CLK_OUT.n585 CLK_OUT.n584 1.1005
R4949 CLK_OUT.n583 CLK_OUT.n363 1.1005
R4950 CLK_OUT.n580 CLK_OUT.n579 1.1005
R4951 CLK_OUT.n576 CLK_OUT.n575 1.1005
R4952 CLK_OUT.n569 CLK_OUT.n369 1.1005
R4953 CLK_OUT.n571 CLK_OUT.n570 1.1005
R4954 CLK_OUT.n568 CLK_OUT.n368 1.1005
R4955 CLK_OUT.n560 CLK_OUT.n374 1.1005
R4956 CLK_OUT.n555 CLK_OUT.n554 1.1005
R4957 CLK_OUT.n553 CLK_OUT.n376 1.1005
R4958 CLK_OUT.n550 CLK_OUT.n377 1.1005
R4959 CLK_OUT.n544 CLK_OUT.n543 1.1005
R4960 CLK_OUT.n540 CLK_OUT.n539 1.1005
R4961 CLK_OUT.n538 CLK_OUT.n381 1.1005
R4962 CLK_OUT.n537 CLK_OUT.n536 1.1005
R4963 CLK_OUT.n384 CLK_OUT.n383 1.1005
R4964 CLK_OUT.n519 CLK_OUT.n388 1.1005
R4965 CLK_OUT.n518 CLK_OUT.n517 1.1005
R4966 CLK_OUT.n390 CLK_OUT.n389 1.1005
R4967 CLK_OUT.n510 CLK_OUT.n509 1.1005
R4968 CLK_OUT.n508 CLK_OUT.n393 1.1005
R4969 CLK_OUT.n507 CLK_OUT.n506 1.1005
R4970 CLK_OUT.n504 CLK_OUT.n503 1.1005
R4971 CLK_OUT.n498 CLK_OUT.n395 1.1005
R4972 CLK_OUT.n495 CLK_OUT.n396 1.1005
R4973 CLK_OUT.n492 CLK_OUT.n397 1.1005
R4974 CLK_OUT.n486 CLK_OUT.n398 1.1005
R4975 CLK_OUT.n485 CLK_OUT.n484 1.1005
R4976 CLK_OUT.n400 CLK_OUT.n399 1.1005
R4977 CLK_OUT.n477 CLK_OUT.n476 1.1005
R4978 CLK_OUT.n475 CLK_OUT.n402 1.1005
R4979 CLK_OUT.n469 CLK_OUT.n403 1.1005
R4980 CLK_OUT.n468 CLK_OUT.n405 1.1005
R4981 CLK_OUT.n467 CLK_OUT.n466 1.1005
R4982 CLK_OUT.n463 CLK_OUT.n462 1.1005
R4983 CLK_OUT.n460 CLK_OUT.n459 1.1005
R4984 CLK_OUT.n453 CLK_OUT.n413 1.1005
R4985 CLK_OUT.n455 CLK_OUT.n454 1.1005
R4986 CLK_OUT.n452 CLK_OUT.n412 1.1005
R4987 CLK_OUT.n447 CLK_OUT.n446 1.1005
R4988 CLK_OUT.n437 CLK_OUT.n417 1.1005
R4989 CLK_OUT.n436 CLK_OUT.n435 1.1005
R4990 CLK_OUT.n427 CLK_OUT.n426 1.1005
R4991 CLK_OUT.n428 CLK_OUT.n427 1.1005
R4992 CLK_OUT.n425 CLK_OUT.n420 1.1005
R4993 CLK_OUT.n419 CLK_OUT.n418 1.1005
R4994 CLK_OUT.n445 CLK_OUT.n415 1.1005
R4995 CLK_OUT.n444 CLK_OUT.n443 1.1005
R4996 CLK_OUT.n442 CLK_OUT.n416 1.1005
R4997 CLK_OUT.n439 CLK_OUT.n438 1.1005
R4998 CLK_OUT.n448 CLK_OUT.n414 1.1005
R4999 CLK_OUT.n451 CLK_OUT.n450 1.1005
R5000 CLK_OUT.n410 CLK_OUT.n409 1.1005
R5001 CLK_OUT.n461 CLK_OUT.n408 1.1005
R5002 CLK_OUT.n407 CLK_OUT.n406 1.1005
R5003 CLK_OUT.n471 CLK_OUT.n470 1.1005
R5004 CLK_OUT.n478 CLK_OUT.n401 1.1005
R5005 CLK_OUT.n480 CLK_OUT.n479 1.1005
R5006 CLK_OUT.n488 CLK_OUT.n487 1.1005
R5007 CLK_OUT.n494 CLK_OUT.n493 1.1005
R5008 CLK_OUT.n497 CLK_OUT.n496 1.1005
R5009 CLK_OUT.n505 CLK_OUT.n394 1.1005
R5010 CLK_OUT.n511 CLK_OUT.n392 1.1005
R5011 CLK_OUT.n513 CLK_OUT.n512 1.1005
R5012 CLK_OUT.n521 CLK_OUT.n520 1.1005
R5013 CLK_OUT.n529 CLK_OUT.n528 1.1005
R5014 CLK_OUT.n527 CLK_OUT.n385 1.1005
R5015 CLK_OUT.n526 CLK_OUT.n525 1.1005
R5016 CLK_OUT.n387 CLK_OUT.n386 1.1005
R5017 CLK_OUT.n534 CLK_OUT.n533 1.1005
R5018 CLK_OUT.n535 CLK_OUT.n382 1.1005
R5019 CLK_OUT.n541 CLK_OUT.n380 1.1005
R5020 CLK_OUT.n542 CLK_OUT.n378 1.1005
R5021 CLK_OUT.n552 CLK_OUT.n551 1.1005
R5022 CLK_OUT.n562 CLK_OUT.n561 1.1005
R5023 CLK_OUT.n559 CLK_OUT.n373 1.1005
R5024 CLK_OUT.n558 CLK_OUT.n557 1.1005
R5025 CLK_OUT.n556 CLK_OUT.n375 1.1005
R5026 CLK_OUT.n371 CLK_OUT.n370 1.1005
R5027 CLK_OUT.n567 CLK_OUT.n566 1.1005
R5028 CLK_OUT.n367 CLK_OUT.n366 1.1005
R5029 CLK_OUT.n577 CLK_OUT.n365 1.1005
R5030 CLK_OUT.n578 CLK_OUT.n364 1.1005
R5031 CLK_OUT.n592 CLK_OUT.n359 1.1005
R5032 CLK_OUT.n587 CLK_OUT.n360 1.1005
R5033 CLK_OUT.n589 CLK_OUT.n588 1.1005
R5034 CLK_OUT.n586 CLK_OUT.n362 1.1005
R5035 CLK_OUT.n595 CLK_OUT.n358 1.1005
R5036 CLK_OUT.n597 CLK_OUT.n596 1.1005
R5037 CLK_OUT.n605 CLK_OUT.n604 1.1005
R5038 CLK_OUT.n611 CLK_OUT.n610 1.1005
R5039 CLK_OUT.n614 CLK_OUT.n613 1.1005
R5040 CLK_OUT.n622 CLK_OUT.n351 1.1005
R5041 CLK_OUT.n628 CLK_OUT.n349 1.1005
R5042 CLK_OUT.n630 CLK_OUT.n629 1.1005
R5043 CLK_OUT.n638 CLK_OUT.n637 1.1005
R5044 CLK_OUT.n646 CLK_OUT.n645 1.1005
R5045 CLK_OUT.n644 CLK_OUT.n342 1.1005
R5046 CLK_OUT.n643 CLK_OUT.n642 1.1005
R5047 CLK_OUT.n344 CLK_OUT.n343 1.1005
R5048 CLK_OUT.n651 CLK_OUT.n650 1.1005
R5049 CLK_OUT.n652 CLK_OUT.n339 1.1005
R5050 CLK_OUT.n658 CLK_OUT.n337 1.1005
R5051 CLK_OUT.n661 CLK_OUT.n660 1.1005
R5052 CLK_OUT.n670 CLK_OUT.n333 1.1005
R5053 CLK_OUT.n678 CLK_OUT.n331 1.1005
R5054 CLK_OUT.n677 CLK_OUT.n676 1.1005
R5055 CLK_OUT.n675 CLK_OUT.n332 1.1005
R5056 CLK_OUT.n672 CLK_OUT.n671 1.1005
R5057 CLK_OUT.n681 CLK_OUT.n330 1.1005
R5058 CLK_OUT.n684 CLK_OUT.n683 1.1005
R5059 CLK_OUT.n326 CLK_OUT.n325 1.1005
R5060 CLK_OUT.n694 CLK_OUT.n324 1.1005
R5061 CLK_OUT.n695 CLK_OUT.n323 1.1005
R5062 CLK_OUT.n703 CLK_OUT.n321 1.1005
R5063 CLK_OUT.n709 CLK_OUT.n318 1.1005
R5064 CLK_OUT.n319 CLK_OUT.n317 1.1005
R5065 CLK_OUT.n706 CLK_OUT.n705 1.1005
R5066 CLK_OUT.n1336 CLK_OUT.n1335 1.1005
R5067 CLK_OUT.n1334 CLK_OUT.n34 1.1005
R5068 CLK_OUT.n1333 CLK_OUT.n34 1.1005
R5069 CLK_OUT.n708 CLK_OUT.n319 1.1005
R5070 CLK_OUT.n707 CLK_OUT.n706 1.1005
R5071 CLK_OUT.n1337 CLK_OUT.n33 1.1005
R5072 CLK_OUT.n862 CLK_OUT.n861 1.1005
R5073 CLK_OUT.n860 CLK_OUT.n274 1.1005
R5074 CLK_OUT.n859 CLK_OUT.n858 1.1005
R5075 CLK_OUT.n279 CLK_OUT.n278 1.1005
R5076 CLK_OUT.n836 CLK_OUT.n280 1.1005
R5077 CLK_OUT.n838 CLK_OUT.n837 1.1005
R5078 CLK_OUT.n835 CLK_OUT.n834 1.1005
R5079 CLK_OUT.n826 CLK_OUT.n283 1.1005
R5080 CLK_OUT.n819 CLK_OUT.n818 1.1005
R5081 CLK_OUT.n817 CLK_OUT.n816 1.1005
R5082 CLK_OUT.n809 CLK_OUT.n287 1.1005
R5083 CLK_OUT.n802 CLK_OUT.n801 1.1005
R5084 CLK_OUT.n800 CLK_OUT.n799 1.1005
R5085 CLK_OUT.n791 CLK_OUT.n291 1.1005
R5086 CLK_OUT.n784 CLK_OUT.n783 1.1005
R5087 CLK_OUT.n782 CLK_OUT.n781 1.1005
R5088 CLK_OUT.n296 CLK_OUT.n295 1.1005
R5089 CLK_OUT.n757 CLK_OUT.n297 1.1005
R5090 CLK_OUT.n758 CLK_OUT.n299 1.1005
R5091 CLK_OUT.n760 CLK_OUT.n759 1.1005
R5092 CLK_OUT.n756 CLK_OUT.n755 1.1005
R5093 CLK_OUT.n745 CLK_OUT.n301 1.1005
R5094 CLK_OUT.n310 CLK_OUT.n304 1.1005
R5095 CLK_OUT.n311 CLK_OUT.n305 1.1005
R5096 CLK_OUT.n312 CLK_OUT.n306 1.1005
R5097 CLK_OUT.n313 CLK_OUT.n308 1.1005
R5098 CLK_OUT.n720 CLK_OUT.n309 1.1005
R5099 CLK_OUT.n717 CLK_OUT.n716 1.1005
R5100 CLK_OUT.n433 CLK_OUT.n432 0.733833
R5101 CLK_OUT.n1185 CLK_OUT.n1184 0.733833
R5102 CLK_OUT.n1338 CLK_OUT.n1337 0.733833
R5103 CLK_OUT.n716 CLK_OUT.n715 0.733833
R5104 CLK_OUT.n1103 CLK_OUT.n126 0.573769
R5105 CLK_OUT.n992 CLK_OUT.n179 0.573769
R5106 CLK_OUT.n139 CLK_OUT.n137 0.573695
R5107 CLK_OUT.n192 CLK_OUT.n190 0.573695
R5108 CLK_OUT.n1051 CLK_OUT.n150 0.573346
R5109 CLK_OUT.n424 CLK_OUT.n420 0.550549
R5110 CLK_OUT.n704 CLK_OUT.n319 0.550549
R5111 CLK_OUT.n1107 CLK_OUT.n125 0.39244
R5112 CLK_OUT.n996 CLK_OUT.n178 0.39244
R5113 CLK_OUT.n1081 CLK_OUT.n138 0.389994
R5114 CLK_OUT.n970 CLK_OUT.n191 0.389994
R5115 CLK_OUT.n1055 CLK_OUT.n149 0.387191
R5116 CLK_OUT.n1143 CLK_OUT.n107 0.384705
R5117 CLK_OUT.n1032 CLK_OUT.n1031 0.384705
R5118 CLK_OUT.n1108 CLK_OUT.n122 0.384705
R5119 CLK_OUT.n997 CLK_OUT.n175 0.384705
R5120 CLK_OUT.n1142 CLK_OUT.n110 0.382331
R5121 CLK_OUT.n1029 CLK_OUT.n162 0.382331
R5122 CLK_OUT.n1115 CLK_OUT.n111 0.382034
R5123 CLK_OUT.n1004 CLK_OUT.n163 0.382034
R5124 CLK_OUT.n1090 CLK_OUT.n127 0.379547
R5125 CLK_OUT.n1045 CLK_OUT.n151 0.379547
R5126 CLK_OUT.n979 CLK_OUT.n180 0.379547
R5127 CLK_OUT.n1059 CLK_OUT.n140 0.376968
R5128 CLK_OUT.n1063 CLK_OUT.n140 0.376876
R5129 CLK_OUT.n1092 CLK_OUT.n127 0.375976
R5130 CLK_OUT.n981 CLK_OUT.n180 0.375976
R5131 CLK_OUT.n154 CLK_OUT.n151 0.375884
R5132 CLK_OUT.n1117 CLK_OUT.n111 0.374982
R5133 CLK_OUT.n1006 CLK_OUT.n163 0.374982
R5134 CLK_OUT.n1142 CLK_OUT.n109 0.374889
R5135 CLK_OUT.n1029 CLK_OUT.n161 0.374889
R5136 CLK_OUT.n1143 CLK_OUT.n108 0.373984
R5137 CLK_OUT.n1031 CLK_OUT.n158 0.373984
R5138 CLK_OUT.n1109 CLK_OUT.n1108 0.373891
R5139 CLK_OUT.n998 CLK_OUT.n997 0.373891
R5140 CLK_OUT CLK_OUT.n1372 0.323045
R5141 CLK_OUT.n1184 CLK_OUT.n1183 0.275034
R5142 CLK_OUT.n1198 CLK_OUT.n74 0.0405
R5143 CLK_OUT.n1198 CLK_OUT.n72 0.0405
R5144 CLK_OUT.n1202 CLK_OUT.n72 0.0405
R5145 CLK_OUT.n1202 CLK_OUT.n62 0.0405
R5146 CLK_OUT.n1218 CLK_OUT.n62 0.0405
R5147 CLK_OUT.n1218 CLK_OUT.n60 0.0405
R5148 CLK_OUT.n1222 CLK_OUT.n60 0.0405
R5149 CLK_OUT.n1222 CLK_OUT.n2 0.0405
R5150 CLK_OUT.n1370 CLK_OUT.n2 0.0405
R5151 CLK_OUT.n1370 CLK_OUT.n1369 0.0405
R5152 CLK_OUT.n1369 CLK_OUT.n1368 0.0405
R5153 CLK_OUT.n1368 CLK_OUT.n6 0.0405
R5154 CLK_OUT.n1364 CLK_OUT.n6 0.0405
R5155 CLK_OUT.n1364 CLK_OUT.n1363 0.0405
R5156 CLK_OUT.n1362 CLK_OUT.n11 0.0405
R5157 CLK_OUT.n1358 CLK_OUT.n11 0.0405
R5158 CLK_OUT.n1358 CLK_OUT.n1357 0.0405
R5159 CLK_OUT.n1357 CLK_OUT.n1356 0.0405
R5160 CLK_OUT.n1356 CLK_OUT.n16 0.0405
R5161 CLK_OUT.n1352 CLK_OUT.n16 0.0405
R5162 CLK_OUT.n1352 CLK_OUT.n1351 0.0405
R5163 CLK_OUT.n1351 CLK_OUT.n1350 0.0405
R5164 CLK_OUT.n1350 CLK_OUT.n21 0.0405
R5165 CLK_OUT.n1346 CLK_OUT.n21 0.0405
R5166 CLK_OUT.n1346 CLK_OUT.n1345 0.0405
R5167 CLK_OUT.n1345 CLK_OUT.n1344 0.0405
R5168 CLK_OUT.n957 CLK_OUT.n956 0.0405
R5169 CLK_OUT.n956 CLK_OUT.n955 0.0405
R5170 CLK_OUT.n955 CLK_OUT.n201 0.0405
R5171 CLK_OUT.n951 CLK_OUT.n201 0.0405
R5172 CLK_OUT.n951 CLK_OUT.n950 0.0405
R5173 CLK_OUT.n950 CLK_OUT.n949 0.0405
R5174 CLK_OUT.n949 CLK_OUT.n206 0.0405
R5175 CLK_OUT.n945 CLK_OUT.n206 0.0405
R5176 CLK_OUT.n945 CLK_OUT.n944 0.0405
R5177 CLK_OUT.n944 CLK_OUT.n943 0.0405
R5178 CLK_OUT.n943 CLK_OUT.n211 0.0405
R5179 CLK_OUT.n939 CLK_OUT.n211 0.0405
R5180 CLK_OUT.n939 CLK_OUT.n938 0.0405
R5181 CLK_OUT.n938 CLK_OUT.n937 0.0405
R5182 CLK_OUT.n933 CLK_OUT.n216 0.0405
R5183 CLK_OUT.n933 CLK_OUT.n932 0.0405
R5184 CLK_OUT.n932 CLK_OUT.n931 0.0405
R5185 CLK_OUT.n931 CLK_OUT.n221 0.0405
R5186 CLK_OUT.n927 CLK_OUT.n221 0.0405
R5187 CLK_OUT.n927 CLK_OUT.n926 0.0405
R5188 CLK_OUT.n926 CLK_OUT.n925 0.0405
R5189 CLK_OUT.n925 CLK_OUT.n226 0.0405
R5190 CLK_OUT.n921 CLK_OUT.n226 0.0405
R5191 CLK_OUT.n921 CLK_OUT.n920 0.0405
R5192 CLK_OUT.n920 CLK_OUT.n919 0.0405
R5193 CLK_OUT.n919 CLK_OUT.n231 0.0405
R5194 CLK_OUT.n958 CLK_OUT.n197 0.0405
R5195 CLK_OUT.n954 CLK_OUT.n197 0.0405
R5196 CLK_OUT.n954 CLK_OUT.n953 0.0405
R5197 CLK_OUT.n953 CLK_OUT.n952 0.0405
R5198 CLK_OUT.n952 CLK_OUT.n202 0.0405
R5199 CLK_OUT.n948 CLK_OUT.n202 0.0405
R5200 CLK_OUT.n948 CLK_OUT.n947 0.0405
R5201 CLK_OUT.n947 CLK_OUT.n946 0.0405
R5202 CLK_OUT.n946 CLK_OUT.n207 0.0405
R5203 CLK_OUT.n942 CLK_OUT.n207 0.0405
R5204 CLK_OUT.n942 CLK_OUT.n941 0.0405
R5205 CLK_OUT.n941 CLK_OUT.n940 0.0405
R5206 CLK_OUT.n940 CLK_OUT.n212 0.0405
R5207 CLK_OUT.n936 CLK_OUT.n212 0.0405
R5208 CLK_OUT.n935 CLK_OUT.n934 0.0405
R5209 CLK_OUT.n934 CLK_OUT.n217 0.0405
R5210 CLK_OUT.n930 CLK_OUT.n217 0.0405
R5211 CLK_OUT.n930 CLK_OUT.n929 0.0405
R5212 CLK_OUT.n929 CLK_OUT.n928 0.0405
R5213 CLK_OUT.n928 CLK_OUT.n222 0.0405
R5214 CLK_OUT.n924 CLK_OUT.n222 0.0405
R5215 CLK_OUT.n924 CLK_OUT.n923 0.0405
R5216 CLK_OUT.n923 CLK_OUT.n922 0.0405
R5217 CLK_OUT.n922 CLK_OUT.n227 0.0405
R5218 CLK_OUT.n918 CLK_OUT.n227 0.0405
R5219 CLK_OUT.n918 CLK_OUT.n917 0.0405
R5220 CLK_OUT.n1199 CLK_OUT.n73 0.0405
R5221 CLK_OUT.n1200 CLK_OUT.n1199 0.0405
R5222 CLK_OUT.n1201 CLK_OUT.n1200 0.0405
R5223 CLK_OUT.n1201 CLK_OUT.n61 0.0405
R5224 CLK_OUT.n1219 CLK_OUT.n61 0.0405
R5225 CLK_OUT.n1220 CLK_OUT.n1219 0.0405
R5226 CLK_OUT.n1221 CLK_OUT.n1220 0.0405
R5227 CLK_OUT.n1221 CLK_OUT.n0 0.0405
R5228 CLK_OUT.n1371 CLK_OUT.n1 0.0405
R5229 CLK_OUT.n1367 CLK_OUT.n1 0.0405
R5230 CLK_OUT.n1367 CLK_OUT.n1366 0.0405
R5231 CLK_OUT.n1366 CLK_OUT.n1365 0.0405
R5232 CLK_OUT.n1365 CLK_OUT.n7 0.0405
R5233 CLK_OUT.n1361 CLK_OUT.n1360 0.0405
R5234 CLK_OUT.n1360 CLK_OUT.n1359 0.0405
R5235 CLK_OUT.n1359 CLK_OUT.n12 0.0405
R5236 CLK_OUT.n1355 CLK_OUT.n12 0.0405
R5237 CLK_OUT.n1355 CLK_OUT.n1354 0.0405
R5238 CLK_OUT.n1354 CLK_OUT.n1353 0.0405
R5239 CLK_OUT.n1353 CLK_OUT.n17 0.0405
R5240 CLK_OUT.n1349 CLK_OUT.n17 0.0405
R5241 CLK_OUT.n1349 CLK_OUT.n1348 0.0405
R5242 CLK_OUT.n1348 CLK_OUT.n1347 0.0405
R5243 CLK_OUT.n1347 CLK_OUT.n22 0.0405
R5244 CLK_OUT.n1343 CLK_OUT.n22 0.0405
R5245 CLK_OUT.n1363 CLK_OUT.n1362 0.0360676
R5246 CLK_OUT.n937 CLK_OUT.n216 0.0360676
R5247 CLK_OUT.n936 CLK_OUT.n935 0.0360676
R5248 CLK_OUT.n961 CLK_OUT.n960 0.0360676
R5249 CLK_OUT.n961 CLK_OUT.n184 0.0360676
R5250 CLK_OUT.n986 CLK_OUT.n184 0.0360676
R5251 CLK_OUT.n987 CLK_OUT.n986 0.0360676
R5252 CLK_OUT.n988 CLK_OUT.n987 0.0360676
R5253 CLK_OUT.n988 CLK_OUT.n171 0.0360676
R5254 CLK_OUT.n1011 CLK_OUT.n171 0.0360676
R5255 CLK_OUT.n1012 CLK_OUT.n1011 0.0360676
R5256 CLK_OUT.n1013 CLK_OUT.n1012 0.0360676
R5257 CLK_OUT.n1014 CLK_OUT.n1013 0.0360676
R5258 CLK_OUT.n1015 CLK_OUT.n1014 0.0360676
R5259 CLK_OUT.n1016 CLK_OUT.n1015 0.0360676
R5260 CLK_OUT.n1017 CLK_OUT.n1016 0.0360676
R5261 CLK_OUT.n1017 CLK_OUT.n144 0.0360676
R5262 CLK_OUT.n1069 CLK_OUT.n144 0.0360676
R5263 CLK_OUT.n1070 CLK_OUT.n1069 0.0360676
R5264 CLK_OUT.n1071 CLK_OUT.n1070 0.0360676
R5265 CLK_OUT.n1072 CLK_OUT.n1071 0.0360676
R5266 CLK_OUT.n1072 CLK_OUT.n131 0.0360676
R5267 CLK_OUT.n1097 CLK_OUT.n131 0.0360676
R5268 CLK_OUT.n1098 CLK_OUT.n1097 0.0360676
R5269 CLK_OUT.n1099 CLK_OUT.n1098 0.0360676
R5270 CLK_OUT.n1099 CLK_OUT.n118 0.0360676
R5271 CLK_OUT.n1122 CLK_OUT.n118 0.0360676
R5272 CLK_OUT.n1123 CLK_OUT.n1122 0.0360676
R5273 CLK_OUT.n1124 CLK_OUT.n1123 0.0360676
R5274 CLK_OUT.n1125 CLK_OUT.n1124 0.0360676
R5275 CLK_OUT.n1126 CLK_OUT.n1125 0.0360676
R5276 CLK_OUT.n1126 CLK_OUT.n96 0.0360676
R5277 CLK_OUT.n1169 CLK_OUT.n96 0.0360676
R5278 CLK_OUT.n1170 CLK_OUT.n1169 0.0360676
R5279 CLK_OUT.n1171 CLK_OUT.n1170 0.0360676
R5280 CLK_OUT.n1173 CLK_OUT.n1171 0.0360676
R5281 CLK_OUT.n963 CLK_OUT.n962 0.0360676
R5282 CLK_OUT.n962 CLK_OUT.n185 0.0360676
R5283 CLK_OUT.n985 CLK_OUT.n185 0.0360676
R5284 CLK_OUT.n985 CLK_OUT.n183 0.0360676
R5285 CLK_OUT.n989 CLK_OUT.n183 0.0360676
R5286 CLK_OUT.n989 CLK_OUT.n172 0.0360676
R5287 CLK_OUT.n1010 CLK_OUT.n172 0.0360676
R5288 CLK_OUT.n1010 CLK_OUT.n170 0.0360676
R5289 CLK_OUT.n1022 CLK_OUT.n170 0.0360676
R5290 CLK_OUT.n1022 CLK_OUT.n1021 0.0360676
R5291 CLK_OUT.n1021 CLK_OUT.n1020 0.0360676
R5292 CLK_OUT.n1020 CLK_OUT.n1019 0.0360676
R5293 CLK_OUT.n1019 CLK_OUT.n1018 0.0360676
R5294 CLK_OUT.n1018 CLK_OUT.n145 0.0360676
R5295 CLK_OUT.n1068 CLK_OUT.n145 0.0360676
R5296 CLK_OUT.n1068 CLK_OUT.n143 0.0360676
R5297 CLK_OUT.n1074 CLK_OUT.n143 0.0360676
R5298 CLK_OUT.n1074 CLK_OUT.n1073 0.0360676
R5299 CLK_OUT.n1073 CLK_OUT.n132 0.0360676
R5300 CLK_OUT.n1096 CLK_OUT.n132 0.0360676
R5301 CLK_OUT.n1096 CLK_OUT.n130 0.0360676
R5302 CLK_OUT.n1100 CLK_OUT.n130 0.0360676
R5303 CLK_OUT.n1100 CLK_OUT.n119 0.0360676
R5304 CLK_OUT.n1121 CLK_OUT.n119 0.0360676
R5305 CLK_OUT.n1121 CLK_OUT.n117 0.0360676
R5306 CLK_OUT.n1135 CLK_OUT.n117 0.0360676
R5307 CLK_OUT.n1135 CLK_OUT.n1134 0.0360676
R5308 CLK_OUT.n1134 CLK_OUT.n1127 0.0360676
R5309 CLK_OUT.n1127 CLK_OUT.n97 0.0360676
R5310 CLK_OUT.n1168 CLK_OUT.n97 0.0360676
R5311 CLK_OUT.n1168 CLK_OUT.n95 0.0360676
R5312 CLK_OUT.n1175 CLK_OUT.n95 0.0360676
R5313 CLK_OUT.n1175 CLK_OUT.n1174 0.0360676
R5314 CLK_OUT.n914 CLK_OUT.n913 0.0360676
R5315 CLK_OUT.n913 CLK_OUT.n912 0.0360676
R5316 CLK_OUT.n912 CLK_OUT.n237 0.0360676
R5317 CLK_OUT.n908 CLK_OUT.n237 0.0360676
R5318 CLK_OUT.n908 CLK_OUT.n907 0.0360676
R5319 CLK_OUT.n907 CLK_OUT.n906 0.0360676
R5320 CLK_OUT.n906 CLK_OUT.n242 0.0360676
R5321 CLK_OUT.n902 CLK_OUT.n242 0.0360676
R5322 CLK_OUT.n902 CLK_OUT.n901 0.0360676
R5323 CLK_OUT.n901 CLK_OUT.n900 0.0360676
R5324 CLK_OUT.n900 CLK_OUT.n247 0.0360676
R5325 CLK_OUT.n896 CLK_OUT.n247 0.0360676
R5326 CLK_OUT.n896 CLK_OUT.n895 0.0360676
R5327 CLK_OUT.n895 CLK_OUT.n894 0.0360676
R5328 CLK_OUT.n894 CLK_OUT.n252 0.0360676
R5329 CLK_OUT.n890 CLK_OUT.n252 0.0360676
R5330 CLK_OUT.n890 CLK_OUT.n889 0.0360676
R5331 CLK_OUT.n889 CLK_OUT.n888 0.0360676
R5332 CLK_OUT.n888 CLK_OUT.n257 0.0360676
R5333 CLK_OUT.n884 CLK_OUT.n257 0.0360676
R5334 CLK_OUT.n884 CLK_OUT.n883 0.0360676
R5335 CLK_OUT.n883 CLK_OUT.n882 0.0360676
R5336 CLK_OUT.n882 CLK_OUT.n262 0.0360676
R5337 CLK_OUT.n878 CLK_OUT.n262 0.0360676
R5338 CLK_OUT.n878 CLK_OUT.n877 0.0360676
R5339 CLK_OUT.n877 CLK_OUT.n876 0.0360676
R5340 CLK_OUT.n876 CLK_OUT.n267 0.0360676
R5341 CLK_OUT.n872 CLK_OUT.n267 0.0360676
R5342 CLK_OUT.n872 CLK_OUT.n871 0.0360676
R5343 CLK_OUT.n871 CLK_OUT.n870 0.0360676
R5344 CLK_OUT.n870 CLK_OUT.n867 0.0360676
R5345 CLK_OUT.n867 CLK_OUT.n28 0.0360676
R5346 CLK_OUT.n1340 CLK_OUT.n28 0.0360676
R5347 CLK_OUT.n915 CLK_OUT.n233 0.0360676
R5348 CLK_OUT.n911 CLK_OUT.n233 0.0360676
R5349 CLK_OUT.n911 CLK_OUT.n910 0.0360676
R5350 CLK_OUT.n910 CLK_OUT.n909 0.0360676
R5351 CLK_OUT.n909 CLK_OUT.n238 0.0360676
R5352 CLK_OUT.n905 CLK_OUT.n238 0.0360676
R5353 CLK_OUT.n905 CLK_OUT.n904 0.0360676
R5354 CLK_OUT.n904 CLK_OUT.n903 0.0360676
R5355 CLK_OUT.n903 CLK_OUT.n243 0.0360676
R5356 CLK_OUT.n899 CLK_OUT.n243 0.0360676
R5357 CLK_OUT.n899 CLK_OUT.n898 0.0360676
R5358 CLK_OUT.n898 CLK_OUT.n897 0.0360676
R5359 CLK_OUT.n897 CLK_OUT.n248 0.0360676
R5360 CLK_OUT.n893 CLK_OUT.n248 0.0360676
R5361 CLK_OUT.n893 CLK_OUT.n892 0.0360676
R5362 CLK_OUT.n892 CLK_OUT.n891 0.0360676
R5363 CLK_OUT.n891 CLK_OUT.n253 0.0360676
R5364 CLK_OUT.n887 CLK_OUT.n253 0.0360676
R5365 CLK_OUT.n887 CLK_OUT.n886 0.0360676
R5366 CLK_OUT.n886 CLK_OUT.n885 0.0360676
R5367 CLK_OUT.n885 CLK_OUT.n258 0.0360676
R5368 CLK_OUT.n881 CLK_OUT.n258 0.0360676
R5369 CLK_OUT.n881 CLK_OUT.n880 0.0360676
R5370 CLK_OUT.n880 CLK_OUT.n879 0.0360676
R5371 CLK_OUT.n879 CLK_OUT.n263 0.0360676
R5372 CLK_OUT.n875 CLK_OUT.n263 0.0360676
R5373 CLK_OUT.n875 CLK_OUT.n874 0.0360676
R5374 CLK_OUT.n874 CLK_OUT.n873 0.0360676
R5375 CLK_OUT.n873 CLK_OUT.n268 0.0360676
R5376 CLK_OUT.n869 CLK_OUT.n268 0.0360676
R5377 CLK_OUT.n869 CLK_OUT.n868 0.0360676
R5378 CLK_OUT.n868 CLK_OUT.n27 0.0360676
R5379 CLK_OUT.n1341 CLK_OUT.n27 0.0360676
R5380 CLK_OUT.n1361 CLK_OUT.n7 0.0360676
R5381 CLK_OUT.n1373 CLK_OUT 0.02602
R5382 CLK_OUT.n88 CLK_OUT.n74 0.0234189
R5383 CLK_OUT.n957 CLK_OUT.n196 0.0234189
R5384 CLK_OUT.n959 CLK_OUT.n958 0.0234189
R5385 CLK_OUT.n1172 CLK_OUT.n73 0.0234189
R5386 CLK_OUT.n1344 CLK_OUT.n26 0.0233108
R5387 CLK_OUT.n232 CLK_OUT.n231 0.0233108
R5388 CLK_OUT.n917 CLK_OUT.n916 0.0233108
R5389 CLK_OUT.n1343 CLK_OUT.n1342 0.0233108
R5390 CLK_OUT.n960 CLK_OUT.n959 0.0227703
R5391 CLK_OUT.n963 CLK_OUT.n196 0.0227703
R5392 CLK_OUT.n914 CLK_OUT.n232 0.0227703
R5393 CLK_OUT.n916 CLK_OUT.n915 0.0227703
R5394 CLK_OUT.n1372 CLK_OUT.n1371 0.0220135
R5395 CLK_OUT.n1372 CLK_OUT.n0 0.0189865
R5396 CLK_OUT.n83 CLK_OUT.n76 0.0188784
R5397 CLK_OUT.n81 CLK_OUT.n71 0.0188784
R5398 CLK_OUT.n1207 CLK_OUT.n1204 0.0188784
R5399 CLK_OUT.n1205 CLK_OUT.n63 0.0188784
R5400 CLK_OUT.n1216 CLK_OUT.n65 0.0188784
R5401 CLK_OUT.n1230 CLK_OUT.n1229 0.0188784
R5402 CLK_OUT.n1233 CLK_OUT.n1232 0.0188784
R5403 CLK_OUT.n1241 CLK_OUT.n1240 0.0188784
R5404 CLK_OUT.n1246 CLK_OUT.n1245 0.0188784
R5405 CLK_OUT.n1249 CLK_OUT.n1248 0.0188784
R5406 CLK_OUT.n1257 CLK_OUT.n1256 0.0188784
R5407 CLK_OUT.n1262 CLK_OUT.n1261 0.0188784
R5408 CLK_OUT.n1266 CLK_OUT.n1265 0.0188784
R5409 CLK_OUT.n1273 CLK_OUT.n47 0.0188784
R5410 CLK_OUT.n1276 CLK_OUT.n1275 0.0188784
R5411 CLK_OUT.n1281 CLK_OUT.n1280 0.0188784
R5412 CLK_OUT.n1284 CLK_OUT.n1283 0.0188784
R5413 CLK_OUT.n1290 CLK_OUT.n43 0.0188784
R5414 CLK_OUT.n1301 CLK_OUT.n1300 0.0188784
R5415 CLK_OUT.n1311 CLK_OUT.n1310 0.0188784
R5416 CLK_OUT.n1315 CLK_OUT.n1314 0.0188784
R5417 CLK_OUT.n1319 CLK_OUT.n1318 0.0188784
R5418 CLK_OUT.n1324 CLK_OUT.n1323 0.0188784
R5419 CLK_OUT.n457 CLK_OUT.n456 0.0188784
R5420 CLK_OUT.n465 CLK_OUT.n464 0.0188784
R5421 CLK_OUT.n474 CLK_OUT.n473 0.0188784
R5422 CLK_OUT.n483 CLK_OUT.n482 0.0188784
R5423 CLK_OUT.n490 CLK_OUT.n489 0.0188784
R5424 CLK_OUT.n516 CLK_OUT.n515 0.0188784
R5425 CLK_OUT.n524 CLK_OUT.n523 0.0188784
R5426 CLK_OUT.n531 CLK_OUT.n530 0.0188784
R5427 CLK_OUT.n546 CLK_OUT.n379 0.0188784
R5428 CLK_OUT.n549 CLK_OUT.n548 0.0188784
R5429 CLK_OUT.n563 CLK_OUT.n372 0.0188784
R5430 CLK_OUT.n573 CLK_OUT.n572 0.0188784
R5431 CLK_OUT.n582 CLK_OUT.n581 0.0188784
R5432 CLK_OUT.n591 CLK_OUT.n590 0.0188784
R5433 CLK_OUT.n600 CLK_OUT.n599 0.0188784
R5434 CLK_OUT.n607 CLK_OUT.n606 0.0188784
R5435 CLK_OUT.n618 CLK_OUT.n616 0.0188784
R5436 CLK_OUT.n632 CLK_OUT.n348 0.0188784
R5437 CLK_OUT.n648 CLK_OUT.n647 0.0188784
R5438 CLK_OUT.n663 CLK_OUT.n336 0.0188784
R5439 CLK_OUT.n666 CLK_OUT.n665 0.0188784
R5440 CLK_OUT.n674 CLK_OUT.n673 0.0188784
R5441 CLK_OUT.n689 CLK_OUT.n327 0.0188784
R5442 CLK_OUT.n433 CLK_OUT.n195 0.0188784
R5443 CLK_OUT.n966 CLK_OUT.n965 0.0188784
R5444 CLK_OUT.n975 CLK_OUT.n974 0.0188784
R5445 CLK_OUT.n977 CLK_OUT.n186 0.0188784
R5446 CLK_OUT.n1061 CLK_OUT.n142 0.0188784
R5447 CLK_OUT.n1077 CLK_OUT.n1076 0.0188784
R5448 CLK_OUT.n1086 CLK_OUT.n1085 0.0188784
R5449 CLK_OUT.n1088 CLK_OUT.n133 0.0188784
R5450 CLK_OUT.n715 CLK_OUT.n714 0.0188784
R5451 CLK_OUT.n724 CLK_OUT.n723 0.0188784
R5452 CLK_OUT.n728 CLK_OUT.n727 0.0188784
R5453 CLK_OUT.n732 CLK_OUT.n307 0.0188784
R5454 CLK_OUT.n793 CLK_OUT.n792 0.0188784
R5455 CLK_OUT.n797 CLK_OUT.n796 0.0188784
R5456 CLK_OUT.n804 CLK_OUT.n289 0.0188784
R5457 CLK_OUT.n807 CLK_OUT.n806 0.0188784
R5458 CLK_OUT.n1188 CLK_OUT.n75 0.0187703
R5459 CLK_OUT.n1196 CLK_OUT.n76 0.0187703
R5460 CLK_OUT.n1224 CLK_OUT.n59 0.0187703
R5461 CLK_OUT.n1229 CLK_OUT.n57 0.0187703
R5462 CLK_OUT.n1258 CLK_OUT.n1257 0.0187703
R5463 CLK_OUT.n1295 CLK_OUT.n43 0.0187703
R5464 CLK_OUT.n1298 CLK_OUT.n1297 0.0187703
R5465 CLK_OUT.n1325 CLK_OUT.n1324 0.0187703
R5466 CLK_OUT.n1329 CLK_OUT.n1328 0.0187703
R5467 CLK_OUT.n441 CLK_OUT.n440 0.0187703
R5468 CLK_OUT.n456 CLK_OUT.n411 0.0187703
R5469 CLK_OUT.n501 CLK_OUT.n499 0.0187703
R5470 CLK_OUT.n515 CLK_OUT.n391 0.0187703
R5471 CLK_OUT.n564 CLK_OUT.n563 0.0187703
R5472 CLK_OUT.n633 CLK_OUT.n632 0.0187703
R5473 CLK_OUT.n641 CLK_OUT.n640 0.0187703
R5474 CLK_OUT.n690 CLK_OUT.n689 0.0187703
R5475 CLK_OUT.n699 CLK_OUT.n698 0.0187703
R5476 CLK_OUT.n991 CLK_OUT.n182 0.0187703
R5477 CLK_OUT.n1000 CLK_OUT.n176 0.0187703
R5478 CLK_OUT.n1002 CLK_OUT.n173 0.0187703
R5479 CLK_OUT.n1008 CLK_OUT.n174 0.0187703
R5480 CLK_OUT.n1025 CLK_OUT.n1024 0.0187703
R5481 CLK_OUT.n169 CLK_OUT.n167 0.0187703
R5482 CLK_OUT.n1035 CLK_OUT.n1034 0.0187703
R5483 CLK_OUT.n1039 CLK_OUT.n1038 0.0187703
R5484 CLK_OUT.n1043 CLK_OUT.n1042 0.0187703
R5485 CLK_OUT.n1048 CLK_OUT.n1047 0.0187703
R5486 CLK_OUT.n1050 CLK_OUT.n146 0.0187703
R5487 CLK_OUT.n1066 CLK_OUT.n147 0.0187703
R5488 CLK_OUT.n1102 CLK_OUT.n129 0.0187703
R5489 CLK_OUT.n1111 CLK_OUT.n123 0.0187703
R5490 CLK_OUT.n1113 CLK_OUT.n120 0.0187703
R5491 CLK_OUT.n1119 CLK_OUT.n121 0.0187703
R5492 CLK_OUT.n1138 CLK_OUT.n1137 0.0187703
R5493 CLK_OUT.n1129 CLK_OUT.n116 0.0187703
R5494 CLK_OUT.n1132 CLK_OUT.n1130 0.0187703
R5495 CLK_OUT.n1148 CLK_OUT.n1147 0.0187703
R5496 CLK_OUT.n1150 CLK_OUT.n98 0.0187703
R5497 CLK_OUT.n1166 CLK_OUT.n99 0.0187703
R5498 CLK_OUT.n1158 CLK_OUT.n94 0.0187703
R5499 CLK_OUT.n1178 CLK_OUT.n1177 0.0187703
R5500 CLK_OUT.n738 CLK_OUT.n737 0.0187703
R5501 CLK_OUT.n742 CLK_OUT.n741 0.0187703
R5502 CLK_OUT.n747 CLK_OUT.n303 0.0187703
R5503 CLK_OUT.n750 CLK_OUT.n749 0.0187703
R5504 CLK_OUT.n753 CLK_OUT.n752 0.0187703
R5505 CLK_OUT.n763 CLK_OUT.n762 0.0187703
R5506 CLK_OUT.n767 CLK_OUT.n766 0.0187703
R5507 CLK_OUT.n771 CLK_OUT.n770 0.0187703
R5508 CLK_OUT.n775 CLK_OUT.n774 0.0187703
R5509 CLK_OUT.n779 CLK_OUT.n778 0.0187703
R5510 CLK_OUT.n786 CLK_OUT.n293 0.0187703
R5511 CLK_OUT.n789 CLK_OUT.n788 0.0187703
R5512 CLK_OUT.n814 CLK_OUT.n813 0.0187703
R5513 CLK_OUT.n821 CLK_OUT.n285 0.0187703
R5514 CLK_OUT.n824 CLK_OUT.n823 0.0187703
R5515 CLK_OUT.n829 CLK_OUT.n828 0.0187703
R5516 CLK_OUT.n832 CLK_OUT.n831 0.0187703
R5517 CLK_OUT.n841 CLK_OUT.n840 0.0187703
R5518 CLK_OUT.n845 CLK_OUT.n844 0.0187703
R5519 CLK_OUT.n849 CLK_OUT.n848 0.0187703
R5520 CLK_OUT.n856 CLK_OUT.n855 0.0187703
R5521 CLK_OUT.n853 CLK_OUT.n272 0.0187703
R5522 CLK_OUT.n865 CLK_OUT.n273 0.0187703
R5523 CLK_OUT.n276 CLK_OUT.n29 0.0187703
R5524 CLK_OUT.n82 CLK_OUT.n81 0.0185541
R5525 CLK_OUT.n1319 CLK_OUT.n23 0.0185541
R5526 CLK_OUT.n464 CLK_OUT.n200 0.0185541
R5527 CLK_OUT.n673 CLK_OUT.n229 0.0185541
R5528 CLK_OUT.n983 CLK_OUT.n187 0.0184459
R5529 CLK_OUT.n1094 CLK_OUT.n134 0.0184459
R5530 CLK_OUT.n734 CLK_OUT.n239 0.0184459
R5531 CLK_OUT.n810 CLK_OUT.n260 0.0184459
R5532 CLK_OUT.n1261 CLK_OUT.n8 0.0182297
R5533 CLK_OUT.n572 CLK_OUT.n214 0.0182297
R5534 CLK_OUT.n984 CLK_OUT.n983 0.0181216
R5535 CLK_OUT.n1095 CLK_OUT.n1094 0.0181216
R5536 CLK_OUT.n734 CLK_OUT.n733 0.0181216
R5537 CLK_OUT.n810 CLK_OUT.n259 0.0181216
R5538 CLK_OUT.n1224 CLK_OUT.n1223 0.0175811
R5539 CLK_OUT.n1297 CLK_OUT.n1296 0.0175811
R5540 CLK_OUT.n501 CLK_OUT.n500 0.0175811
R5541 CLK_OUT.n640 CLK_OUT.n223 0.0175811
R5542 CLK_OUT.n991 CLK_OUT.n990 0.0173649
R5543 CLK_OUT.n1102 CLK_OUT.n1101 0.0173649
R5544 CLK_OUT.n738 CLK_OUT.n240 0.0173649
R5545 CLK_OUT.n814 CLK_OUT.n261 0.0173649
R5546 CLK_OUT CLK_OUT.n1374 0.0171486
R5547 CLK_OUT.n977 CLK_OUT.n976 0.0170405
R5548 CLK_OUT.n1088 CLK_OUT.n1087 0.0170405
R5549 CLK_OUT.n307 CLK_OUT.n236 0.0170405
R5550 CLK_OUT.n806 CLK_OUT.n805 0.0170405
R5551 CLK_OUT.n1233 CLK_OUT.n1231 0.0167162
R5552 CLK_OUT.n1283 CLK_OUT.n15 0.0167162
R5553 CLK_OUT.n523 CLK_OUT.n208 0.0167162
R5554 CLK_OUT.n618 CLK_OUT.n617 0.0167162
R5555 CLK_OUT.n1001 CLK_OUT.n1000 0.0162838
R5556 CLK_OUT.n1112 CLK_OUT.n1111 0.0162838
R5557 CLK_OUT.n742 CLK_OUT.n241 0.0162838
R5558 CLK_OUT.n822 CLK_OUT.n821 0.0162838
R5559 CLK_OUT.n1248 CLK_OUT.n51 0.0159595
R5560 CLK_OUT.n47 CLK_OUT.n10 0.0159595
R5561 CLK_OUT.n548 CLK_OUT.n213 0.0159595
R5562 CLK_OUT.n590 CLK_OUT.n361 0.0159595
R5563 CLK_OUT.n974 CLK_OUT.n189 0.0159595
R5564 CLK_OUT.n1085 CLK_OUT.n136 0.0159595
R5565 CLK_OUT.n727 CLK_OUT.n235 0.0159595
R5566 CLK_OUT.n289 CLK_OUT.n256 0.0159595
R5567 CLK_OUT.n1197 CLK_OUT.n75 0.0157432
R5568 CLK_OUT.n1328 CLK_OUT.n24 0.0157432
R5569 CLK_OUT.n440 CLK_OUT.n199 0.0157432
R5570 CLK_OUT.n698 CLK_OUT.n230 0.0157432
R5571 CLK_OUT.n1204 CLK_OUT.n1203 0.0152027
R5572 CLK_OUT.n1315 CLK_OUT.n38 0.0152027
R5573 CLK_OUT.n473 CLK_OUT.n404 0.0152027
R5574 CLK_OUT.n665 CLK_OUT.n228 0.0152027
R5575 CLK_OUT.n1009 CLK_OUT.n173 0.0152027
R5576 CLK_OUT.n1120 CLK_OUT.n120 0.0152027
R5577 CLK_OUT.n748 CLK_OUT.n747 0.0152027
R5578 CLK_OUT.n824 CLK_OUT.n264 0.0152027
R5579 CLK_OUT.n1265 CLK_OUT.n9 0.0148784
R5580 CLK_OUT.n581 CLK_OUT.n215 0.0148784
R5581 CLK_OUT.n965 CLK_OUT.n964 0.0148784
R5582 CLK_OUT.n1076 CLK_OUT.n1075 0.0148784
R5583 CLK_OUT.n723 CLK_OUT.n234 0.0148784
R5584 CLK_OUT.n796 CLK_OUT.n255 0.0148784
R5585 CLK_OUT.n65 CLK_OUT.n64 0.0141216
R5586 CLK_OUT.n1301 CLK_OUT.n18 0.0141216
R5587 CLK_OUT.n489 CLK_OUT.n205 0.0141216
R5588 CLK_OUT.n647 CLK_OUT.n224 0.0141216
R5589 CLK_OUT.n174 CLK_OUT.n166 0.0141216
R5590 CLK_OUT.n121 CLK_OUT.n114 0.0141216
R5591 CLK_OUT.n750 CLK_OUT.n244 0.0141216
R5592 CLK_OUT.n829 CLK_OUT.n265 0.0141216
R5593 CLK_OUT.n1173 CLK_OUT.n1172 0.0137973
R5594 CLK_OUT.n1174 CLK_OUT.n88 0.0137973
R5595 CLK_OUT.n1061 CLK_OUT.n1060 0.0137973
R5596 CLK_OUT.n1185 CLK_OUT.n87 0.0137973
R5597 CLK_OUT.n792 CLK_OUT.n254 0.0137973
R5598 CLK_OUT.n1339 CLK_OUT.n1338 0.0137973
R5599 CLK_OUT.n1340 CLK_OUT.n26 0.0137973
R5600 CLK_OUT.n1342 CLK_OUT.n1341 0.0137973
R5601 CLK_OUT.n861 CLK_OUT.n33 0.0134381
R5602 CLK_OUT.n1240 CLK_OUT.n3 0.0133649
R5603 CLK_OUT.n1281 CLK_OUT.n14 0.0133649
R5604 CLK_OUT.n530 CLK_OUT.n209 0.0133649
R5605 CLK_OUT.n606 CLK_OUT.n220 0.0133649
R5606 CLK_OUT.n1024 CLK_OUT.n1023 0.0130405
R5607 CLK_OUT.n1137 CLK_OUT.n1136 0.0130405
R5608 CLK_OUT.n752 CLK_OUT.n245 0.0130405
R5609 CLK_OUT.n831 CLK_OUT.n266 0.0130405
R5610 CLK_OUT.n1067 CLK_OUT.n1066 0.0128243
R5611 CLK_OUT.n1178 CLK_OUT.n1176 0.0128243
R5612 CLK_OUT.n788 CLK_OUT.n787 0.0128243
R5613 CLK_OUT.n276 CLK_OUT.n275 0.0128243
R5614 CLK_OUT.n1246 CLK_OUT.n5 0.0126081
R5615 CLK_OUT.n1275 CLK_OUT.n1274 0.0126081
R5616 CLK_OUT.n547 CLK_OUT.n546 0.0126081
R5617 CLK_OUT.n599 CLK_OUT.n218 0.0126081
R5618 CLK_OUT.n1187 CLK_OUT.n1186 0.0123919
R5619 CLK_OUT.n30 CLK_OUT.n25 0.0123919
R5620 CLK_OUT.n434 CLK_OUT.n198 0.0123919
R5621 CLK_OUT.n712 CLK_OUT.n320 0.0123919
R5622 CLK_OUT.n167 CLK_OUT.n159 0.0119595
R5623 CLK_OUT.n1133 CLK_OUT.n1129 0.0119595
R5624 CLK_OUT.n763 CLK_OUT.n246 0.0119595
R5625 CLK_OUT.n841 CLK_OUT.n281 0.0119595
R5626 CLK_OUT.n1206 CLK_OUT.n1205 0.0118514
R5627 CLK_OUT.n1311 CLK_OUT.n20 0.0118514
R5628 CLK_OUT.n482 CLK_OUT.n203 0.0118514
R5629 CLK_OUT.n664 CLK_OUT.n663 0.0118514
R5630 CLK_OUT.n1050 CLK_OUT.n1049 0.0117432
R5631 CLK_OUT.n1158 CLK_OUT.n1157 0.0117432
R5632 CLK_OUT.n293 CLK_OUT.n251 0.0117432
R5633 CLK_OUT.n866 CLK_OUT.n865 0.0117432
R5634 CLK_OUT.n1183 CLK_OUT.n85 0.0116588
R5635 CLK_OUT.n1186 CLK_OUT.n1185 0.011527
R5636 CLK_OUT.n434 CLK_OUT.n433 0.011527
R5637 CLK_OUT.n1338 CLK_OUT.n30 0.0114189
R5638 CLK_OUT.n715 CLK_OUT.n712 0.0114189
R5639 CLK_OUT.n313 CLK_OUT.n312 0.0109762
R5640 CLK_OUT.n311 CLK_OUT.n310 0.0109762
R5641 CLK_OUT.n756 CLK_OUT.n301 0.0109762
R5642 CLK_OUT.n759 CLK_OUT.n758 0.0109762
R5643 CLK_OUT.n757 CLK_OUT.n295 0.0109762
R5644 CLK_OUT.n783 CLK_OUT.n782 0.0109762
R5645 CLK_OUT.n800 CLK_OUT.n291 0.0109762
R5646 CLK_OUT.n801 CLK_OUT.n287 0.0109762
R5647 CLK_OUT.n818 CLK_OUT.n817 0.0109762
R5648 CLK_OUT.n835 CLK_OUT.n283 0.0109762
R5649 CLK_OUT.n837 CLK_OUT.n836 0.0109762
R5650 CLK_OUT.n859 CLK_OUT.n278 0.0109762
R5651 CLK_OUT.n861 CLK_OUT.n860 0.0109762
R5652 CLK_OUT.n1192 CLK_OUT.n1191 0.0109762
R5653 CLK_OUT.n1192 CLK_OUT.n67 0.0109762
R5654 CLK_OUT.n1210 CLK_OUT.n67 0.0109762
R5655 CLK_OUT.n1211 CLK_OUT.n1210 0.0109762
R5656 CLK_OUT.n1212 CLK_OUT.n1211 0.0109762
R5657 CLK_OUT.n1212 CLK_OUT.n55 0.0109762
R5658 CLK_OUT.n1236 CLK_OUT.n55 0.0109762
R5659 CLK_OUT.n1237 CLK_OUT.n1236 0.0109762
R5660 CLK_OUT.n1237 CLK_OUT.n53 0.0109762
R5661 CLK_OUT.n1252 CLK_OUT.n53 0.0109762
R5662 CLK_OUT.n1253 CLK_OUT.n1252 0.0109762
R5663 CLK_OUT.n1269 CLK_OUT.n49 0.0109762
R5664 CLK_OUT.n1270 CLK_OUT.n1269 0.0109762
R5665 CLK_OUT.n1270 CLK_OUT.n45 0.0109762
R5666 CLK_OUT.n1287 CLK_OUT.n45 0.0109762
R5667 CLK_OUT.n1288 CLK_OUT.n1287 0.0109762
R5668 CLK_OUT.n1288 CLK_OUT.n41 0.0109762
R5669 CLK_OUT.n1304 CLK_OUT.n41 0.0109762
R5670 CLK_OUT.n1307 CLK_OUT.n1304 0.0109762
R5671 CLK_OUT.n1307 CLK_OUT.n1306 0.0109762
R5672 CLK_OUT.n1306 CLK_OUT.n1305 0.0109762
R5673 CLK_OUT.n1305 CLK_OUT.n35 0.0109762
R5674 CLK_OUT.n1332 CLK_OUT.n35 0.0109762
R5675 CLK_OUT.n971 CLK_OUT.n180 0.0109762
R5676 CLK_OUT.n997 CLK_OUT.n996 0.0109762
R5677 CLK_OUT.n1028 CLK_OUT.n163 0.0109762
R5678 CLK_OUT.n1031 CLK_OUT.n1029 0.0109762
R5679 CLK_OUT.n1030 CLK_OUT.n151 0.0109762
R5680 CLK_OUT.n1056 CLK_OUT.n1055 0.0109762
R5681 CLK_OUT.n1081 CLK_OUT.n140 0.0109762
R5682 CLK_OUT.n1082 CLK_OUT.n127 0.0109762
R5683 CLK_OUT.n1108 CLK_OUT.n1107 0.0109762
R5684 CLK_OUT.n1141 CLK_OUT.n111 0.0109762
R5685 CLK_OUT.n1143 CLK_OUT.n1142 0.0109762
R5686 CLK_OUT.n312 CLK_OUT.n311 0.01095
R5687 CLK_OUT.n310 CLK_OUT.n301 0.01095
R5688 CLK_OUT.n759 CLK_OUT.n756 0.01095
R5689 CLK_OUT.n758 CLK_OUT.n757 0.01095
R5690 CLK_OUT.n782 CLK_OUT.n295 0.01095
R5691 CLK_OUT.n783 CLK_OUT.n291 0.01095
R5692 CLK_OUT.n801 CLK_OUT.n800 0.01095
R5693 CLK_OUT.n817 CLK_OUT.n287 0.01095
R5694 CLK_OUT.n818 CLK_OUT.n283 0.01095
R5695 CLK_OUT.n837 CLK_OUT.n835 0.01095
R5696 CLK_OUT.n836 CLK_OUT.n278 0.01095
R5697 CLK_OUT.n860 CLK_OUT.n859 0.01095
R5698 CLK_OUT.n1253 CLK_OUT.n49 0.01095
R5699 CLK_OUT.n1333 CLK_OUT.n1332 0.01095
R5700 CLK_OUT.n971 CLK_OUT.n970 0.01095
R5701 CLK_OUT.n996 CLK_OUT.n180 0.01095
R5702 CLK_OUT.n997 CLK_OUT.n163 0.01095
R5703 CLK_OUT.n1029 CLK_OUT.n1028 0.01095
R5704 CLK_OUT.n1031 CLK_OUT.n1030 0.01095
R5705 CLK_OUT.n1055 CLK_OUT.n151 0.01095
R5706 CLK_OUT.n1056 CLK_OUT.n140 0.01095
R5707 CLK_OUT.n1082 CLK_OUT.n1081 0.01095
R5708 CLK_OUT.n1107 CLK_OUT.n127 0.01095
R5709 CLK_OUT.n1108 CLK_OUT.n111 0.01095
R5710 CLK_OUT.n1142 CLK_OUT.n1141 0.01095
R5711 CLK_OUT.n1144 CLK_OUT.n1143 0.01095
R5712 CLK_OUT.n1035 CLK_OUT.n157 0.0108784
R5713 CLK_OUT.n1130 CLK_OUT.n105 0.0108784
R5714 CLK_OUT.n767 CLK_OUT.n298 0.0108784
R5715 CLK_OUT.n845 CLK_OUT.n269 0.0108784
R5716 CLK_OUT.n1217 CLK_OUT.n63 0.0107703
R5717 CLK_OUT.n1310 CLK_OUT.n19 0.0107703
R5718 CLK_OUT.n483 CLK_OUT.n204 0.0107703
R5719 CLK_OUT.n336 CLK_OUT.n225 0.0107703
R5720 CLK_OUT.n1047 CLK_OUT.n153 0.0106622
R5721 CLK_OUT.n1167 CLK_OUT.n1166 0.0106622
R5722 CLK_OUT.n778 CLK_OUT.n250 0.0106622
R5723 CLK_OUT.n853 CLK_OUT.n271 0.0106622
R5724 CLK_OUT.n1191 CLK_OUT.n85 0.0106095
R5725 CLK_OUT.n1245 CLK_OUT.n4 0.0100135
R5726 CLK_OUT.n1276 CLK_OUT.n13 0.0100135
R5727 CLK_OUT.n379 CLK_OUT.n210 0.0100135
R5728 CLK_OUT.n600 CLK_OUT.n219 0.0100135
R5729 CLK_OUT.n1039 CLK_OUT.n155 0.0097973
R5730 CLK_OUT.n1149 CLK_OUT.n1148 0.0097973
R5731 CLK_OUT.n771 CLK_OUT.n249 0.0097973
R5732 CLK_OUT.n849 CLK_OUT.n270 0.0097973
R5733 CLK_OUT.n1183 CLK_OUT.n1182 0.00967266
R5734 CLK_OUT.n1042 CLK_OUT.n155 0.00958108
R5735 CLK_OUT.n1150 CLK_OUT.n1149 0.00958108
R5736 CLK_OUT.n774 CLK_OUT.n249 0.00958108
R5737 CLK_OUT.n855 CLK_OUT.n270 0.00958108
R5738 CLK_OUT.n1241 CLK_OUT.n4 0.00925676
R5739 CLK_OUT.n1280 CLK_OUT.n13 0.00925676
R5740 CLK_OUT.n531 CLK_OUT.n210 0.00925676
R5741 CLK_OUT.n607 CLK_OUT.n219 0.00925676
R5742 CLK_OUT.n1055 CLK_OUT.n150 0.00880612
R5743 CLK_OUT.n1043 CLK_OUT.n153 0.00871622
R5744 CLK_OUT.n1167 CLK_OUT.n98 0.00871622
R5745 CLK_OUT.n775 CLK_OUT.n250 0.00871622
R5746 CLK_OUT.n856 CLK_OUT.n271 0.00871622
R5747 CLK_OUT.n1217 CLK_OUT.n1216 0.0085
R5748 CLK_OUT.n1300 CLK_OUT.n19 0.0085
R5749 CLK_OUT.n490 CLK_OUT.n204 0.0085
R5750 CLK_OUT.n648 CLK_OUT.n225 0.0085
R5751 CLK_OUT.n1038 CLK_OUT.n157 0.0085
R5752 CLK_OUT.n1147 CLK_OUT.n105 0.0085
R5753 CLK_OUT.n770 CLK_OUT.n298 0.0085
R5754 CLK_OUT.n848 CLK_OUT.n269 0.0085
R5755 CLK_OUT.n314 CLK_OUT.n313 0.00809524
R5756 CLK_OUT.n1181 CLK_OUT.n91 0.00778095
R5757 CLK_OUT.n1049 CLK_OUT.n1048 0.00763514
R5758 CLK_OUT.n1157 CLK_OUT.n99 0.00763514
R5759 CLK_OUT.n779 CLK_OUT.n251 0.00763514
R5760 CLK_OUT.n866 CLK_OUT.n272 0.00763514
R5761 CLK_OUT.n1207 CLK_OUT.n1206 0.00741892
R5762 CLK_OUT.n1314 CLK_OUT.n20 0.00741892
R5763 CLK_OUT.n474 CLK_OUT.n203 0.00741892
R5764 CLK_OUT.n666 CLK_OUT.n664 0.00741892
R5765 CLK_OUT.n1034 CLK_OUT.n159 0.00741892
R5766 CLK_OUT.n1133 CLK_OUT.n1132 0.00741892
R5767 CLK_OUT.n766 CLK_OUT.n246 0.00741892
R5768 CLK_OUT.n844 CLK_OUT.n281 0.00741892
R5769 CLK_OUT.n1144 CLK_OUT.n103 0.00725714
R5770 CLK_OUT.n1182 CLK_OUT.n1181 0.00707381
R5771 CLK_OUT.n1188 CLK_OUT.n1187 0.00698649
R5772 CLK_OUT.n1329 CLK_OUT.n25 0.00698649
R5773 CLK_OUT.n441 CLK_OUT.n198 0.00698649
R5774 CLK_OUT.n699 CLK_OUT.n320 0.00698649
R5775 CLK_OUT.n970 CLK_OUT.n193 0.00696162
R5776 CLK_OUT.n1335 CLK_OUT.n1333 0.00691667
R5777 CLK_OUT.n1249 CLK_OUT.n5 0.00666216
R5778 CLK_OUT.n1274 CLK_OUT.n1273 0.00666216
R5779 CLK_OUT.n549 CLK_OUT.n547 0.00666216
R5780 CLK_OUT.n591 CLK_OUT.n218 0.00666216
R5781 CLK_OUT.n1067 CLK_OUT.n146 0.00655405
R5782 CLK_OUT.n1176 CLK_OUT.n94 0.00655405
R5783 CLK_OUT.n787 CLK_OUT.n786 0.00655405
R5784 CLK_OUT.n275 CLK_OUT.n273 0.00655405
R5785 CLK_OUT.n1023 CLK_OUT.n169 0.00633784
R5786 CLK_OUT.n1136 CLK_OUT.n116 0.00633784
R5787 CLK_OUT.n762 CLK_OUT.n245 0.00633784
R5788 CLK_OUT.n840 CLK_OUT.n266 0.00633784
R5789 CLK_OUT.n1232 CLK_OUT.n3 0.00590541
R5790 CLK_OUT.n1284 CLK_OUT.n14 0.00590541
R5791 CLK_OUT.n524 CLK_OUT.n209 0.00590541
R5792 CLK_OUT.n616 CLK_OUT.n220 0.00590541
R5793 CLK_OUT.n1081 CLK_OUT.n139 0.00588776
R5794 CLK_OUT.n970 CLK_OUT.n192 0.00588776
R5795 CLK_OUT.n1060 CLK_OUT.n147 0.00547297
R5796 CLK_OUT.n1177 CLK_OUT.n87 0.00547297
R5797 CLK_OUT.n789 CLK_OUT.n254 0.00547297
R5798 CLK_OUT.n1339 CLK_OUT.n29 0.00547297
R5799 CLK_OUT.n1025 CLK_OUT.n166 0.00525676
R5800 CLK_OUT.n1138 CLK_OUT.n114 0.00525676
R5801 CLK_OUT.n753 CLK_OUT.n244 0.00525676
R5802 CLK_OUT.n832 CLK_OUT.n265 0.00525676
R5803 CLK_OUT.n64 CLK_OUT.n59 0.00514865
R5804 CLK_OUT.n1298 CLK_OUT.n18 0.00514865
R5805 CLK_OUT.n499 CLK_OUT.n205 0.00514865
R5806 CLK_OUT.n641 CLK_OUT.n224 0.00514865
R5807 CLK_OUT.n1334 CLK_OUT.n33 0.00440238
R5808 CLK_OUT.n1262 CLK_OUT.n9 0.00439189
R5809 CLK_OUT.n573 CLK_OUT.n215 0.00439189
R5810 CLK_OUT.n964 CLK_OUT.n195 0.00439189
R5811 CLK_OUT.n1075 CLK_OUT.n142 0.00439189
R5812 CLK_OUT.n714 CLK_OUT.n234 0.00439189
R5813 CLK_OUT.n793 CLK_OUT.n255 0.00439189
R5814 CLK_OUT.n1189 CLK_OUT.n86 0.00425921
R5815 CLK_OUT.n1195 CLK_OUT.n77 0.00425921
R5816 CLK_OUT.n70 CLK_OUT.n69 0.00425921
R5817 CLK_OUT.n1215 CLK_OUT.n1214 0.00425921
R5818 CLK_OUT.n1228 CLK_OUT.n56 0.00425921
R5819 CLK_OUT.n1234 CLK_OUT.n54 0.00425921
R5820 CLK_OUT.n1242 CLK_OUT.n1239 0.00425921
R5821 CLK_OUT.n1247 CLK_OUT.n1244 0.00425921
R5822 CLK_OUT.n1263 CLK_OUT.n1260 0.00425921
R5823 CLK_OUT.n1277 CLK_OUT.n46 0.00425921
R5824 CLK_OUT.n1282 CLK_OUT.n1279 0.00425921
R5825 CLK_OUT.n1285 CLK_OUT.n44 0.00425921
R5826 CLK_OUT.n1292 CLK_OUT.n1291 0.00425921
R5827 CLK_OUT.n1302 CLK_OUT.n40 0.00425921
R5828 CLK_OUT.n1312 CLK_OUT.n1309 0.00425921
R5829 CLK_OUT.n1327 CLK_OUT.n1326 0.00425921
R5830 CLK_OUT.n1330 CLK_OUT.n31 0.00425921
R5831 CLK_OUT.n1037 CLK_OUT.n1036 0.00425921
R5832 CLK_OUT.n1041 CLK_OUT.n1040 0.00425921
R5833 CLK_OUT.n1146 CLK_OUT.n106 0.00425921
R5834 CLK_OUT.n1151 CLK_OUT.n104 0.00425921
R5835 CLK_OUT.n731 CLK_OUT.n730 0.00425921
R5836 CLK_OUT.n736 CLK_OUT.n735 0.00425921
R5837 CLK_OUT.n740 CLK_OUT.n739 0.00425921
R5838 CLK_OUT.n744 CLK_OUT.n743 0.00425921
R5839 CLK_OUT.n765 CLK_OUT.n764 0.00425921
R5840 CLK_OUT.n769 CLK_OUT.n768 0.00425921
R5841 CLK_OUT.n773 CLK_OUT.n772 0.00425921
R5842 CLK_OUT.n777 CLK_OUT.n776 0.00425921
R5843 CLK_OUT.n794 CLK_OUT.n791 0.00425921
R5844 CLK_OUT.n808 CLK_OUT.n288 0.00425921
R5845 CLK_OUT.n812 CLK_OUT.n811 0.00425921
R5846 CLK_OUT.n815 CLK_OUT.n286 0.00425921
R5847 CLK_OUT.n820 CLK_OUT.n284 0.00425921
R5848 CLK_OUT.n843 CLK_OUT.n842 0.00425921
R5849 CLK_OUT.n847 CLK_OUT.n846 0.00425921
R5850 CLK_OUT.n851 CLK_OUT.n850 0.00425921
R5851 CLK_OUT.n857 CLK_OUT.n854 0.00425921
R5852 CLK_OUT.n1156 CLK_OUT.n1155 0.00424524
R5853 CLK_OUT.n1195 CLK_OUT.n1194 0.0042371
R5854 CLK_OUT.n84 CLK_OUT.n80 0.0042371
R5855 CLK_OUT.n78 CLK_OUT.n68 0.0042371
R5856 CLK_OUT.n1208 CLK_OUT.n70 0.0042371
R5857 CLK_OUT.n1225 CLK_OUT.n58 0.0042371
R5858 CLK_OUT.n1228 CLK_OUT.n1227 0.0042371
R5859 CLK_OUT.n1250 CLK_OUT.n1247 0.0042371
R5860 CLK_OUT.n1255 CLK_OUT.n52 0.0042371
R5861 CLK_OUT.n1259 CLK_OUT.n50 0.0042371
R5862 CLK_OUT.n1260 CLK_OUT.n1259 0.0042371
R5863 CLK_OUT.n1264 CLK_OUT.n1263 0.0042371
R5864 CLK_OUT.n1267 CLK_OUT.n48 0.0042371
R5865 CLK_OUT.n1272 CLK_OUT.n46 0.0042371
R5866 CLK_OUT.n1294 CLK_OUT.n1292 0.0042371
R5867 CLK_OUT.n1299 CLK_OUT.n42 0.0042371
R5868 CLK_OUT.n1313 CLK_OUT.n1312 0.0042371
R5869 CLK_OUT.n1317 CLK_OUT.n1316 0.0042371
R5870 CLK_OUT.n1322 CLK_OUT.n1320 0.0042371
R5871 CLK_OUT.n1326 CLK_OUT.n36 0.0042371
R5872 CLK_OUT.n978 CLK_OUT.n188 0.0042371
R5873 CLK_OUT.n1007 CLK_OUT.n164 0.0042371
R5874 CLK_OUT.n1026 CLK_OUT.n165 0.0042371
R5875 CLK_OUT.n1065 CLK_OUT.n1064 0.0042371
R5876 CLK_OUT.n1089 CLK_OUT.n135 0.0042371
R5877 CLK_OUT.n1118 CLK_OUT.n112 0.0042371
R5878 CLK_OUT.n1139 CLK_OUT.n113 0.0042371
R5879 CLK_OUT.n1159 CLK_OUT.n92 0.0042371
R5880 CLK_OUT.n1179 CLK_OUT.n93 0.0042371
R5881 CLK_OUT.n726 CLK_OUT.n725 0.0042371
R5882 CLK_OUT.n730 CLK_OUT.n729 0.0042371
R5883 CLK_OUT.n746 CLK_OUT.n744 0.0042371
R5884 CLK_OUT.n751 CLK_OUT.n302 0.0042371
R5885 CLK_OUT.n754 CLK_OUT.n300 0.0042371
R5886 CLK_OUT.n764 CLK_OUT.n761 0.0042371
R5887 CLK_OUT.n780 CLK_OUT.n777 0.0042371
R5888 CLK_OUT.n785 CLK_OUT.n294 0.0042371
R5889 CLK_OUT.n790 CLK_OUT.n292 0.0042371
R5890 CLK_OUT.n791 CLK_OUT.n790 0.0042371
R5891 CLK_OUT.n795 CLK_OUT.n794 0.0042371
R5892 CLK_OUT.n798 CLK_OUT.n290 0.0042371
R5893 CLK_OUT.n803 CLK_OUT.n288 0.0042371
R5894 CLK_OUT.n825 CLK_OUT.n284 0.0042371
R5895 CLK_OUT.n830 CLK_OUT.n827 0.0042371
R5896 CLK_OUT.n833 CLK_OUT.n282 0.0042371
R5897 CLK_OUT.n842 CLK_OUT.n839 0.0042371
R5898 CLK_OUT.n854 CLK_OUT.n852 0.0042371
R5899 CLK_OUT.n864 CLK_OUT.n863 0.0042371
R5900 CLK_OUT.n277 CLK_OUT.n32 0.0042371
R5901 CLK_OUT.n1337 CLK_OUT.n32 0.0042371
R5902 CLK_OUT.n718 CLK_OUT.n717 0.00423273
R5903 CLK_OUT.n429 CLK_OUT.n428 0.00422178
R5904 CLK_OUT.n705 CLK_OUT.n317 0.00422178
R5905 CLK_OUT.n1154 CLK_OUT.n103 0.00421905
R5906 CLK_OUT.n1009 CLK_OUT.n1008 0.00417568
R5907 CLK_OUT.n1120 CLK_OUT.n1119 0.00417568
R5908 CLK_OUT.n749 CLK_OUT.n748 0.00417568
R5909 CLK_OUT.n828 CLK_OUT.n264 0.00417568
R5910 CLK_OUT.n1193 CLK_OUT.n84 0.00410442
R5911 CLK_OUT.n1322 CLK_OUT.n1321 0.00410442
R5912 CLK_OUT.n1203 CLK_OUT.n71 0.00406757
R5913 CLK_OUT.n1318 CLK_OUT.n38 0.00406757
R5914 CLK_OUT.n465 CLK_OUT.n404 0.00406757
R5915 CLK_OUT.n674 CLK_OUT.n228 0.00406757
R5916 CLK_OUT.n1051 CLK_OUT.n148 0.00402269
R5917 CLK_OUT.n982 CLK_OUT.n178 0.00398793
R5918 CLK_OUT.n1093 CLK_OUT.n125 0.00398793
R5919 CLK_OUT.n735 CLK_OUT.n306 0.00397174
R5920 CLK_OUT.n773 CLK_OUT.n296 0.00397174
R5921 CLK_OUT.n811 CLK_OUT.n809 0.00397174
R5922 CLK_OUT.n858 CLK_OUT.n851 0.00397174
R5923 CLK_OUT.n1243 CLK_OUT.n1242 0.00394963
R5924 CLK_OUT.n1279 CLK_OUT.n1278 0.00394963
R5925 CLK_OUT.n973 CLK_OUT.n190 0.00394626
R5926 CLK_OUT.n1084 CLK_OUT.n137 0.00394626
R5927 CLK_OUT.n421 CLK_OUT.n191 0.00393696
R5928 CLK_OUT.n1058 CLK_OUT.n138 0.00393696
R5929 CLK_OUT.n992 CLK_OUT.n177 0.00390294
R5930 CLK_OUT.n1103 CLK_OUT.n124 0.00390294
R5931 CLK_OUT.n1046 CLK_OUT.n149 0.00389381
R5932 CLK_OUT.n1003 CLK_OUT.n175 0.00385851
R5933 CLK_OUT.n1032 CLK_OUT.n160 0.00385851
R5934 CLK_OUT.n1114 CLK_OUT.n122 0.00385851
R5935 CLK_OUT.n1128 CLK_OUT.n107 0.00385851
R5936 CLK_OUT.n1004 CLK_OUT.n1003 0.00380768
R5937 CLK_OUT.n1115 CLK_OUT.n1114 0.00380768
R5938 CLK_OUT.n162 CLK_OUT.n160 0.00380053
R5939 CLK_OUT.n1128 CLK_OUT.n110 0.00380053
R5940 CLK_OUT.n1215 CLK_OUT.n66 0.00379484
R5941 CLK_OUT.n1308 CLK_OUT.n40 0.00379484
R5942 CLK_OUT.n716 CLK_OUT.n316 0.00379484
R5943 CLK_OUT.n1184 CLK_OUT.n90 0.00377273
R5944 CLK_OUT.n979 CLK_OUT.n978 0.0037725
R5945 CLK_OUT.n1046 CLK_OUT.n1045 0.0037725
R5946 CLK_OUT.n1090 CLK_OUT.n1089 0.0037725
R5947 CLK_OUT.n1163 CLK_OUT.n1162 0.00374762
R5948 CLK_OUT.n1059 CLK_OUT.n1058 0.00372958
R5949 CLK_OUT.n745 CLK_OUT.n302 0.0037285
R5950 CLK_OUT.n827 CLK_OUT.n826 0.0037285
R5951 CLK_OUT.n1064 CLK_OUT.n1063 0.00372177
R5952 CLK_OUT.n760 CLK_OUT.n300 0.00370639
R5953 CLK_OUT.n838 CLK_OUT.n282 0.00370639
R5954 CLK_OUT.n1161 CLK_OUT.n91 0.00369524
R5955 CLK_OUT.n1226 CLK_OUT.n1225 0.00366216
R5956 CLK_OUT.n1293 CLK_OUT.n42 0.00366216
R5957 CLK_OUT.n102 CLK_OUT.n100 0.00366216
R5958 CLK_OUT.n1153 CLK_OUT.n1152 0.00364005
R5959 CLK_OUT.n1197 CLK_OUT.n1196 0.00363514
R5960 CLK_OUT.n1325 CLK_OUT.n24 0.00363514
R5961 CLK_OUT.n411 CLK_OUT.n199 0.00363514
R5962 CLK_OUT.n690 CLK_OUT.n230 0.00363514
R5963 CLK_OUT.n721 CLK_OUT.n719 0.00359048
R5964 CLK_OUT.n1041 CLK_OUT.n154 0.00358532
R5965 CLK_OUT.n428 CLK_OUT.n424 0.00357902
R5966 CLK_OUT.n705 CLK_OUT.n704 0.00357902
R5967 CLK_OUT.n982 CLK_OUT.n981 0.00357098
R5968 CLK_OUT.n1093 CLK_OUT.n1092 0.00357098
R5969 CLK_OUT.n1235 CLK_OUT.n1234 0.00348526
R5970 CLK_OUT.n1289 CLK_OUT.n44 0.00348526
R5971 CLK_OUT.n1007 CLK_OUT.n1006 0.003457
R5972 CLK_OUT.n1118 CLK_OUT.n1117 0.003457
R5973 CLK_OUT.n165 CLK_OUT.n161 0.00344926
R5974 CLK_OUT.n113 CLK_OUT.n109 0.00344926
R5975 CLK_OUT.n740 CLK_OUT.n304 0.00344103
R5976 CLK_OUT.n768 CLK_OUT.n299 0.00344103
R5977 CLK_OUT.n819 CLK_OUT.n286 0.00344103
R5978 CLK_OUT.n846 CLK_OUT.n280 0.00344103
R5979 CLK_OUT.n1033 CLK_OUT.n158 0.00343273
R5980 CLK_OUT.n1131 CLK_OUT.n108 0.00343273
R5981 CLK_OUT.n999 CLK_OUT.n998 0.00341839
R5982 CLK_OUT.n1110 CLK_OUT.n1109 0.00341839
R5983 CLK_OUT.n1107 CLK_OUT.n126 0.00341837
R5984 CLK_OUT.n996 CLK_OUT.n179 0.00341837
R5985 CLK_OUT.n720 CLK_OUT.n314 0.00335476
R5986 CLK_OUT.n1209 CLK_OUT.n68 0.00335258
R5987 CLK_OUT.n1316 CLK_OUT.n39 0.00335258
R5988 CLK_OUT.n998 CLK_OUT.n177 0.0033136
R5989 CLK_OUT.n1109 CLK_OUT.n124 0.0033136
R5990 CLK_OUT.n1256 CLK_OUT.n51 0.00331081
R5991 CLK_OUT.n1266 CLK_OUT.n10 0.00331081
R5992 CLK_OUT.n372 CLK_OUT.n213 0.00331081
R5993 CLK_OUT.n582 CLK_OUT.n361 0.00331081
R5994 CLK_OUT.n966 CLK_OUT.n189 0.00331081
R5995 CLK_OUT.n1077 CLK_OUT.n136 0.00331081
R5996 CLK_OUT.n724 CLK_OUT.n235 0.00331081
R5997 CLK_OUT.n797 CLK_OUT.n256 0.00331081
R5998 CLK_OUT.n168 CLK_OUT.n161 0.00330444
R5999 CLK_OUT.n115 CLK_OUT.n109 0.00330444
R6000 CLK_OUT.n1036 CLK_OUT.n158 0.0032992
R6001 CLK_OUT.n108 CLK_OUT.n106 0.0032992
R6002 CLK_OUT.n1006 CLK_OUT.n1005 0.00329663
R6003 CLK_OUT.n1117 CLK_OUT.n1116 0.00329663
R6004 CLK_OUT.n1164 CLK_OUT.n101 0.00324201
R6005 CLK_OUT.n1251 CLK_OUT.n52 0.00319779
R6006 CLK_OUT.n1271 CLK_OUT.n48 0.00319779
R6007 CLK_OUT.n1160 CLK_OUT.n1159 0.00319779
R6008 CLK_OUT.n781 CLK_OUT.n294 0.00319779
R6009 CLK_OUT.n864 CLK_OUT.n274 0.00319779
R6010 CLK_OUT.n973 CLK_OUT.n972 0.00317568
R6011 CLK_OUT.n1084 CLK_OUT.n1083 0.00317568
R6012 CLK_OUT.n726 CLK_OUT.n308 0.00317568
R6013 CLK_OUT.n802 CLK_OUT.n290 0.00317568
R6014 CLK_OUT.n981 CLK_OUT.n980 0.00316007
R6015 CLK_OUT.n1092 CLK_OUT.n1091 0.00316007
R6016 CLK_OUT.n1044 CLK_OUT.n154 0.00314581
R6017 CLK_OUT.n722 CLK_OUT.n315 0.00310934
R6018 CLK_OUT.n1002 CLK_OUT.n1001 0.00309459
R6019 CLK_OUT.n1113 CLK_OUT.n1112 0.00309459
R6020 CLK_OUT.n303 CLK_OUT.n241 0.00309459
R6021 CLK_OUT.n823 CLK_OUT.n822 0.00309459
R6022 CLK_OUT.n1190 CLK_OUT.n1189 0.003043
R6023 CLK_OUT.n1331 CLK_OUT.n1330 0.003043
R6024 CLK_OUT.n1062 CLK_OUT.n1059 0.00302306
R6025 CLK_OUT.n1063 CLK_OUT.n1062 0.00300884
R6026 CLK_OUT.n470 CLK_OUT.n468 0.0029881
R6027 CLK_OUT.n505 CLK_OUT.n504 0.0029881
R6028 CLK_OUT.n520 CLK_OUT.n386 0.0029881
R6029 CLK_OUT.n622 CLK_OUT.n621 0.0029881
R6030 CLK_OUT.n1045 CLK_OUT.n1044 0.00298054
R6031 CLK_OUT.n980 CLK_OUT.n979 0.00298054
R6032 CLK_OUT.n1091 CLK_OUT.n1090 0.00298054
R6033 CLK_OUT.n637 CLK_OUT.n343 0.0029619
R6034 CLK_OUT.n671 CLK_OUT.n670 0.0029619
R6035 CLK_OUT.n168 CLK_OUT.n162 0.00293083
R6036 CLK_OUT.n115 CLK_OUT.n110 0.00293083
R6037 CLK_OUT.n1005 CLK_OUT.n1004 0.0029237
R6038 CLK_OUT.n1116 CLK_OUT.n1115 0.0029237
R6039 CLK_OUT.n1255 CLK_OUT.n1254 0.00291032
R6040 CLK_OUT.n1268 CLK_OUT.n1267 0.00291032
R6041 CLK_OUT.n1057 CLK_OUT.n148 0.00291032
R6042 CLK_OUT.n1180 CLK_OUT.n92 0.00291032
R6043 CLK_OUT.n725 CLK_OUT.n309 0.00291032
R6044 CLK_OUT.n785 CLK_OUT.n784 0.00291032
R6045 CLK_OUT.n799 CLK_OUT.n798 0.00291032
R6046 CLK_OUT.n863 CLK_OUT.n862 0.00291032
R6047 CLK_OUT.n999 CLK_OUT.n175 0.00289527
R6048 CLK_OUT.n1110 CLK_OUT.n122 0.00289527
R6049 CLK_OUT.n1033 CLK_OUT.n1032 0.00289527
R6050 CLK_OUT.n1131 CLK_OUT.n107 0.00289527
R6051 CLK_OUT.n426 CLK_OUT.n424 0.00287188
R6052 CLK_OUT.n707 CLK_OUT.n704 0.00284569
R6053 CLK_OUT.n152 CLK_OUT.n149 0.00283826
R6054 CLK_OUT.n1335 CLK_OUT.n1334 0.00283095
R6055 CLK_OUT.n194 CLK_OUT.n191 0.00279542
R6056 CLK_OUT.n141 CLK_OUT.n138 0.00279542
R6057 CLK_OUT.n181 CLK_OUT.n178 0.00276679
R6058 CLK_OUT.n128 CLK_OUT.n125 0.00276679
R6059 CLK_OUT.n79 CLK_OUT.n78 0.00275553
R6060 CLK_OUT.n1317 CLK_OUT.n37 0.00275553
R6061 CLK_OUT.n89 CLK_OUT.n86 0.00273342
R6062 CLK_OUT.n1337 CLK_OUT.n31 0.00273342
R6063 CLK_OUT.n426 CLK_OUT.n425 0.00272619
R6064 CLK_OUT.n425 CLK_OUT.n418 0.00272619
R6065 CLK_OUT.n444 CLK_OUT.n416 0.00272619
R6066 CLK_OUT.n446 CLK_OUT.n445 0.00272619
R6067 CLK_OUT.n454 CLK_OUT.n453 0.00272619
R6068 CLK_OUT.n462 CLK_OUT.n406 0.00272619
R6069 CLK_OUT.n467 CLK_OUT.n406 0.00272619
R6070 CLK_OUT.n469 CLK_OUT.n402 0.00272619
R6071 CLK_OUT.n477 CLK_OUT.n402 0.00272619
R6072 CLK_OUT.n485 CLK_OUT.n399 0.00272619
R6073 CLK_OUT.n486 CLK_OUT.n485 0.00272619
R6074 CLK_OUT.n495 CLK_OUT.n494 0.00272619
R6075 CLK_OUT.n496 CLK_OUT.n495 0.00272619
R6076 CLK_OUT.n506 CLK_OUT.n393 0.00272619
R6077 CLK_OUT.n510 CLK_OUT.n393 0.00272619
R6078 CLK_OUT.n518 CLK_OUT.n389 0.00272619
R6079 CLK_OUT.n519 CLK_OUT.n518 0.00272619
R6080 CLK_OUT.n527 CLK_OUT.n526 0.00272619
R6081 CLK_OUT.n528 CLK_OUT.n383 0.00272619
R6082 CLK_OUT.n540 CLK_OUT.n381 0.00272619
R6083 CLK_OUT.n552 CLK_OUT.n377 0.00272619
R6084 CLK_OUT.n553 CLK_OUT.n552 0.00272619
R6085 CLK_OUT.n559 CLK_OUT.n558 0.00272619
R6086 CLK_OUT.n561 CLK_OUT.n559 0.00272619
R6087 CLK_OUT.n561 CLK_OUT.n560 0.00272619
R6088 CLK_OUT.n570 CLK_OUT.n569 0.00272619
R6089 CLK_OUT.n579 CLK_OUT.n578 0.00272619
R6090 CLK_OUT.n578 CLK_OUT.n363 0.00272619
R6091 CLK_OUT.n588 CLK_OUT.n587 0.00272619
R6092 CLK_OUT.n587 CLK_OUT.n359 0.00272619
R6093 CLK_OUT.n594 CLK_OUT.n359 0.00272619
R6094 CLK_OUT.n602 CLK_OUT.n356 0.00272619
R6095 CLK_OUT.n603 CLK_OUT.n602 0.00272619
R6096 CLK_OUT.n612 CLK_OUT.n611 0.00272619
R6097 CLK_OUT.n613 CLK_OUT.n612 0.00272619
R6098 CLK_OUT.n627 CLK_OUT.n350 0.00272619
R6099 CLK_OUT.n636 CLK_OUT.n635 0.00272619
R6100 CLK_OUT.n644 CLK_OUT.n643 0.00272619
R6101 CLK_OUT.n645 CLK_OUT.n340 0.00272619
R6102 CLK_OUT.n657 CLK_OUT.n338 0.00272619
R6103 CLK_OUT.n669 CLK_OUT.n334 0.00272619
R6104 CLK_OUT.n670 CLK_OUT.n669 0.00272619
R6105 CLK_OUT.n677 CLK_OUT.n332 0.00272619
R6106 CLK_OUT.n678 CLK_OUT.n677 0.00272619
R6107 CLK_OUT.n679 CLK_OUT.n678 0.00272619
R6108 CLK_OUT.n687 CLK_OUT.n685 0.00272619
R6109 CLK_OUT.n687 CLK_OUT.n686 0.00272619
R6110 CLK_OUT.n696 CLK_OUT.n694 0.00272619
R6111 CLK_OUT.n696 CLK_OUT.n695 0.00272619
R6112 CLK_OUT.n710 CLK_OUT.n709 0.00272619
R6113 CLK_OUT.n708 CLK_OUT.n707 0.00272619
R6114 CLK_OUT.n436 CLK_OUT.n418 0.0027
R6115 CLK_OUT.n445 CLK_OUT.n444 0.0027
R6116 CLK_OUT.n454 CLK_OUT.n452 0.0027
R6117 CLK_OUT.n462 CLK_OUT.n461 0.0027
R6118 CLK_OUT.n470 CLK_OUT.n469 0.0027
R6119 CLK_OUT.n496 CLK_OUT.n395 0.0027
R6120 CLK_OUT.n528 CLK_OUT.n527 0.0027
R6121 CLK_OUT.n536 CLK_OUT.n381 0.0027
R6122 CLK_OUT.n542 CLK_OUT.n377 0.0027
R6123 CLK_OUT.n570 CLK_OUT.n568 0.0027
R6124 CLK_OUT.n579 CLK_OUT.n577 0.0027
R6125 CLK_OUT.n613 CLK_OUT.n352 0.0027
R6126 CLK_OUT.n623 CLK_OUT.n350 0.0027
R6127 CLK_OUT.n635 CLK_OUT.n346 0.0027
R6128 CLK_OUT.n645 CLK_OUT.n644 0.0027
R6129 CLK_OUT.n653 CLK_OUT.n338 0.0027
R6130 CLK_OUT.n659 CLK_OUT.n334 0.0027
R6131 CLK_OUT.n695 CLK_OUT.n322 0.0027
R6132 CLK_OUT.n709 CLK_OUT.n708 0.0027
R6133 CLK_OUT.n504 CLK_OUT.n395 0.00264762
R6134 CLK_OUT.n643 CLK_OUT.n343 0.00264762
R6135 CLK_OUT.n739 CLK_OUT.n305 0.00264496
R6136 CLK_OUT.n816 CLK_OUT.n815 0.00264496
R6137 CLK_OUT.n1037 CLK_OUT.n156 0.00262285
R6138 CLK_OUT.n1146 CLK_OUT.n1145 0.00262285
R6139 CLK_OUT.n769 CLK_OUT.n297 0.00262285
R6140 CLK_OUT.n847 CLK_OUT.n279 0.00262285
R6141 CLK_OUT.n520 CLK_OUT.n519 0.00262143
R6142 CLK_OUT.n623 CLK_OUT.n622 0.00262143
R6143 CLK_OUT.n1238 CLK_OUT.n54 0.00260074
R6144 CLK_OUT.n1286 CLK_OUT.n1285 0.00260074
R6145 CLK_OUT.n472 CLK_OUT.n405 0.00257862
R6146 CLK_OUT.n672 CLK_OUT.n333 0.00257862
R6147 CLK_OUT.n621 CLK_OUT.n352 0.00256905
R6148 CLK_OUT.n1231 CLK_OUT.n1230 0.00255405
R6149 CLK_OUT.n1290 CLK_OUT.n15 0.00255405
R6150 CLK_OUT.n516 CLK_OUT.n208 0.00255405
R6151 CLK_OUT.n617 CLK_OUT.n348 0.00255405
R6152 CLK_OUT.n526 CLK_OUT.n386 0.00254286
R6153 CLK_OUT.n637 CLK_OUT.n636 0.00254286
R6154 CLK_OUT.n522 CLK_OUT.n387 0.0025344
R6155 CLK_OUT.n506 CLK_OUT.n505 0.00251667
R6156 CLK_OUT.n620 CLK_OUT.n619 0.00251228
R6157 CLK_OUT.n431 CLK_OUT.n430 0.0024936
R6158 CLK_OUT.n468 CLK_OUT.n467 0.00246429
R6159 CLK_OUT.n671 CLK_OUT.n332 0.00246429
R6160 CLK_OUT.n1213 CLK_OUT.n58 0.00244595
R6161 CLK_OUT.n1303 CLK_OUT.n1299 0.00244595
R6162 CLK_OUT.n487 CLK_OUT.n486 0.0024381
R6163 CLK_OUT.n653 CLK_OUT.n652 0.0024381
R6164 CLK_OUT.n503 CLK_OUT.n502 0.00242383
R6165 CLK_OUT.n639 CLK_OUT.n344 0.00242383
R6166 CLK_OUT.n719 CLK_OUT.n718 0.00238571
R6167 CLK_OUT.n1163 CLK_OUT.n1156 0.00238571
R6168 CLK_OUT.n451 CLK_OUT.n414 0.00238571
R6169 CLK_OUT.n460 CLK_OUT.n409 0.00238571
R6170 CLK_OUT.n479 CLK_OUT.n478 0.00238571
R6171 CLK_OUT.n487 CLK_OUT.n397 0.00238571
R6172 CLK_OUT.n512 CLK_OUT.n511 0.00238571
R6173 CLK_OUT.n535 CLK_OUT.n534 0.00238571
R6174 CLK_OUT.n543 CLK_OUT.n541 0.00238571
R6175 CLK_OUT.n567 CLK_OUT.n370 0.00238571
R6176 CLK_OUT.n576 CLK_OUT.n366 0.00238571
R6177 CLK_OUT.n585 CLK_OUT.n363 0.00238571
R6178 CLK_OUT.n596 CLK_OUT.n595 0.00238571
R6179 CLK_OUT.n604 CLK_OUT.n354 0.00238571
R6180 CLK_OUT.n629 CLK_OUT.n628 0.00238571
R6181 CLK_OUT.n652 CLK_OUT.n651 0.00238571
R6182 CLK_OUT.n660 CLK_OUT.n658 0.00238571
R6183 CLK_OUT.n684 CLK_OUT.n330 0.00238571
R6184 CLK_OUT.n693 CLK_OUT.n325 0.00238571
R6185 CLK_OUT.n443 CLK_OUT.n442 0.00237961
R6186 CLK_OUT.n447 CLK_OUT.n415 0.00237961
R6187 CLK_OUT.n455 CLK_OUT.n413 0.00237961
R6188 CLK_OUT.n463 CLK_OUT.n407 0.00237961
R6189 CLK_OUT.n466 CLK_OUT.n407 0.00237961
R6190 CLK_OUT.n475 CLK_OUT.n403 0.00237961
R6191 CLK_OUT.n476 CLK_OUT.n475 0.00237961
R6192 CLK_OUT.n484 CLK_OUT.n400 0.00237961
R6193 CLK_OUT.n484 CLK_OUT.n398 0.00237961
R6194 CLK_OUT.n493 CLK_OUT.n396 0.00237961
R6195 CLK_OUT.n497 CLK_OUT.n396 0.00237961
R6196 CLK_OUT.n508 CLK_OUT.n507 0.00237961
R6197 CLK_OUT.n509 CLK_OUT.n508 0.00237961
R6198 CLK_OUT.n517 CLK_OUT.n390 0.00237961
R6199 CLK_OUT.n517 CLK_OUT.n388 0.00237961
R6200 CLK_OUT.n525 CLK_OUT.n385 0.00237961
R6201 CLK_OUT.n529 CLK_OUT.n384 0.00237961
R6202 CLK_OUT.n539 CLK_OUT.n538 0.00237961
R6203 CLK_OUT.n551 CLK_OUT.n550 0.00237961
R6204 CLK_OUT.n551 CLK_OUT.n376 0.00237961
R6205 CLK_OUT.n557 CLK_OUT.n373 0.00237961
R6206 CLK_OUT.n562 CLK_OUT.n373 0.00237961
R6207 CLK_OUT.n562 CLK_OUT.n374 0.00237961
R6208 CLK_OUT.n571 CLK_OUT.n369 0.00237961
R6209 CLK_OUT.n580 CLK_OUT.n364 0.00237961
R6210 CLK_OUT.n583 CLK_OUT.n364 0.00237961
R6211 CLK_OUT.n589 CLK_OUT.n360 0.00237961
R6212 CLK_OUT.n592 CLK_OUT.n360 0.00237961
R6213 CLK_OUT.n593 CLK_OUT.n592 0.00237961
R6214 CLK_OUT.n601 CLK_OUT.n357 0.00237961
R6215 CLK_OUT.n601 CLK_OUT.n355 0.00237961
R6216 CLK_OUT.n610 CLK_OUT.n353 0.00237961
R6217 CLK_OUT.n614 CLK_OUT.n353 0.00237961
R6218 CLK_OUT.n626 CLK_OUT.n625 0.00237961
R6219 CLK_OUT.n634 CLK_OUT.n345 0.00237961
R6220 CLK_OUT.n642 CLK_OUT.n342 0.00237961
R6221 CLK_OUT.n646 CLK_OUT.n341 0.00237961
R6222 CLK_OUT.n656 CLK_OUT.n655 0.00237961
R6223 CLK_OUT.n668 CLK_OUT.n667 0.00237961
R6224 CLK_OUT.n668 CLK_OUT.n333 0.00237961
R6225 CLK_OUT.n676 CLK_OUT.n675 0.00237961
R6226 CLK_OUT.n676 CLK_OUT.n331 0.00237961
R6227 CLK_OUT.n680 CLK_OUT.n331 0.00237961
R6228 CLK_OUT.n688 CLK_OUT.n328 0.00237961
R6229 CLK_OUT.n688 CLK_OUT.n329 0.00237961
R6230 CLK_OUT.n697 CLK_OUT.n324 0.00237961
R6231 CLK_OUT.n697 CLK_OUT.n323 0.00237961
R6232 CLK_OUT.n711 CLK_OUT.n318 0.00237961
R6233 CLK_OUT.n432 CLK_OUT.n423 0.00237961
R6234 CLK_OUT.n968 CLK_OUT.n967 0.00237961
R6235 CLK_OUT.n1027 CLK_OUT.n164 0.00237961
R6236 CLK_OUT.n1027 CLK_OUT.n1026 0.00237961
R6237 CLK_OUT.n1053 CLK_OUT.n1052 0.00237961
R6238 CLK_OUT.n1079 CLK_OUT.n1078 0.00237961
R6239 CLK_OUT.n1140 CLK_OUT.n112 0.00237961
R6240 CLK_OUT.n1140 CLK_OUT.n1139 0.00237961
R6241 CLK_OUT.n755 CLK_OUT.n751 0.00237961
R6242 CLK_OUT.n755 CLK_OUT.n754 0.00237961
R6243 CLK_OUT.n834 CLK_OUT.n830 0.00237961
R6244 CLK_OUT.n834 CLK_OUT.n833 0.00237961
R6245 CLK_OUT.n536 CLK_OUT.n535 0.00235952
R6246 CLK_OUT.n558 CLK_OUT.n375 0.00235952
R6247 CLK_OUT.n435 CLK_OUT.n419 0.00235749
R6248 CLK_OUT.n443 CLK_OUT.n415 0.00235749
R6249 CLK_OUT.n455 CLK_OUT.n412 0.00235749
R6250 CLK_OUT.n463 CLK_OUT.n408 0.00235749
R6251 CLK_OUT.n471 CLK_OUT.n403 0.00235749
R6252 CLK_OUT.n498 CLK_OUT.n497 0.00235749
R6253 CLK_OUT.n529 CLK_OUT.n385 0.00235749
R6254 CLK_OUT.n538 CLK_OUT.n537 0.00235749
R6255 CLK_OUT.n550 CLK_OUT.n378 0.00235749
R6256 CLK_OUT.n571 CLK_OUT.n368 0.00235749
R6257 CLK_OUT.n580 CLK_OUT.n365 0.00235749
R6258 CLK_OUT.n615 CLK_OUT.n614 0.00235749
R6259 CLK_OUT.n625 CLK_OUT.n624 0.00235749
R6260 CLK_OUT.n634 CLK_OUT.n347 0.00235749
R6261 CLK_OUT.n646 CLK_OUT.n342 0.00235749
R6262 CLK_OUT.n655 CLK_OUT.n654 0.00235749
R6263 CLK_OUT.n667 CLK_OUT.n335 0.00235749
R6264 CLK_OUT.n700 CLK_OUT.n323 0.00235749
R6265 CLK_OUT.n994 CLK_OUT.n993 0.00235749
R6266 CLK_OUT.n1105 CLK_OUT.n1104 0.00235749
R6267 CLK_OUT.n604 CLK_OUT.n603 0.00233333
R6268 CLK_OUT.n503 CLK_OUT.n498 0.00231327
R6269 CLK_OUT.n642 CLK_OUT.n344 0.00231327
R6270 CLK_OUT.n437 CLK_OUT.n436 0.00230714
R6271 CLK_OUT.n702 CLK_OUT.n322 0.00230714
R6272 CLK_OUT.n710 CLK_OUT.n703 0.00230714
R6273 CLK_OUT.n1214 CLK_OUT.n1213 0.00229115
R6274 CLK_OUT.n1303 CLK_OUT.n1302 0.00229115
R6275 CLK_OUT.n521 CLK_OUT.n388 0.00229115
R6276 CLK_OUT.n624 CLK_OUT.n351 0.00229115
R6277 CLK_OUT.n438 CLK_OUT.n416 0.00228095
R6278 CLK_OUT.n453 CLK_OUT.n409 0.00228095
R6279 CLK_OUT.n685 CLK_OUT.n684 0.00225476
R6280 CLK_OUT.n620 CLK_OUT.n615 0.00224693
R6281 CLK_OUT.n976 CLK_OUT.n975 0.00222973
R6282 CLK_OUT.n1087 CLK_OUT.n1086 0.00222973
R6283 CLK_OUT.n728 CLK_OUT.n236 0.00222973
R6284 CLK_OUT.n805 CLK_OUT.n804 0.00222973
R6285 CLK_OUT.n525 CLK_OUT.n387 0.00222482
R6286 CLK_OUT.n638 CLK_OUT.n345 0.00222482
R6287 CLK_OUT.n507 CLK_OUT.n394 0.0022027
R6288 CLK_OUT.n554 CLK_OUT.n553 0.00220238
R6289 CLK_OUT.n588 CLK_OUT.n586 0.00220238
R6290 CLK_OUT.n568 CLK_OUT.n567 0.00217619
R6291 CLK_OUT.n569 CLK_OUT.n366 0.00217619
R6292 CLK_OUT.n466 CLK_OUT.n405 0.00215848
R6293 CLK_OUT.n675 CLK_OUT.n672 0.00215848
R6294 CLK_OUT.n1239 CLK_OUT.n1238 0.00213636
R6295 CLK_OUT.n1286 CLK_OUT.n1282 0.00213636
R6296 CLK_OUT.n488 CLK_OUT.n398 0.00213636
R6297 CLK_OUT.n654 CLK_OUT.n339 0.00213636
R6298 CLK_OUT.n1040 CLK_OUT.n156 0.00211425
R6299 CLK_OUT.n1145 CLK_OUT.n104 0.00211425
R6300 CLK_OUT.n772 CLK_OUT.n297 0.00211425
R6301 CLK_OUT.n850 CLK_OUT.n279 0.00211425
R6302 CLK_OUT.n721 CLK_OUT.n720 0.00209762
R6303 CLK_OUT.n452 CLK_OUT.n451 0.00209762
R6304 CLK_OUT.n584 CLK_OUT.n583 0.00209214
R6305 CLK_OUT.n995 CLK_OUT.n181 0.00209214
R6306 CLK_OUT.n1106 CLK_OUT.n128 0.00209214
R6307 CLK_OUT.n736 CLK_OUT.n305 0.00209214
R6308 CLK_OUT.n816 CLK_OUT.n812 0.00209214
R6309 CLK_OUT.n686 CLK_OUT.n325 0.00207143
R6310 CLK_OUT.n537 CLK_OUT.n382 0.00207002
R6311 CLK_OUT.n557 CLK_OUT.n556 0.00207002
R6312 CLK_OUT.n605 CLK_OUT.n355 0.00204791
R6313 CLK_OUT.n435 CLK_OUT.n417 0.0020258
R6314 CLK_OUT.n701 CLK_OUT.n700 0.0020258
R6315 CLK_OUT.n711 CLK_OUT.n321 0.0020258
R6316 CLK_OUT.n541 CLK_OUT.n540 0.00201905
R6317 CLK_OUT.n990 CLK_OUT.n176 0.00201351
R6318 CLK_OUT.n1101 CLK_OUT.n123 0.00201351
R6319 CLK_OUT.n741 CLK_OUT.n240 0.00201351
R6320 CLK_OUT.n285 CLK_OUT.n261 0.00201351
R6321 CLK_OUT.n80 CLK_OUT.n79 0.00200369
R6322 CLK_OUT.n1320 CLK_OUT.n37 0.00200369
R6323 CLK_OUT.n442 CLK_OUT.n439 0.00200369
R6324 CLK_OUT.n413 CLK_OUT.n410 0.00200369
R6325 CLK_OUT.n431 CLK_OUT.n429 0.00200107
R6326 CLK_OUT.n430 CLK_OUT.n193 0.00200107
R6327 CLK_OUT.n717 CLK_OUT.n317 0.00200107
R6328 CLK_OUT.n596 CLK_OUT.n356 0.00199286
R6329 CLK_OUT.n683 CLK_OUT.n328 0.00198157
R6330 CLK_OUT.n555 CLK_OUT.n376 0.00193735
R6331 CLK_OUT.n589 CLK_OUT.n362 0.00193735
R6332 CLK_OUT.n566 CLK_OUT.n368 0.00191523
R6333 CLK_OUT.n369 CLK_OUT.n367 0.00191523
R6334 CLK_OUT.n432 CLK_OUT.n420 0.00191523
R6335 CLK_OUT.n423 CLK_OUT.n422 0.00191523
R6336 CLK_OUT.n716 CLK_OUT.n319 0.00191523
R6337 CLK_OUT.n1337 CLK_OUT.n1336 0.00191523
R6338 CLK_OUT.n479 CLK_OUT.n399 0.00191429
R6339 CLK_OUT.n658 CLK_OUT.n657 0.00191429
R6340 CLK_OUT.n492 CLK_OUT.n491 0.00187101
R6341 CLK_OUT.n993 CLK_OUT.n992 0.00185493
R6342 CLK_OUT.n1104 CLK_OUT.n1103 0.00185493
R6343 CLK_OUT.n1254 CLK_OUT.n50 0.00184889
R6344 CLK_OUT.n1268 CLK_OUT.n1264 0.00184889
R6345 CLK_OUT.n450 CLK_OUT.n412 0.00184889
R6346 CLK_OUT.n650 CLK_OUT.n649 0.00184889
R6347 CLK_OUT.n969 CLK_OUT.n194 0.00184889
R6348 CLK_OUT.n1065 CLK_OUT.n1057 0.00184889
R6349 CLK_OUT.n1080 CLK_OUT.n141 0.00184889
R6350 CLK_OUT.n1180 CLK_OUT.n1179 0.00184889
R6351 CLK_OUT.n722 CLK_OUT.n309 0.00184889
R6352 CLK_OUT.n784 CLK_OUT.n292 0.00184889
R6353 CLK_OUT.n799 CLK_OUT.n795 0.00184889
R6354 CLK_OUT.n862 CLK_OUT.n277 0.00184889
R6355 CLK_OUT.n629 CLK_OUT.n346 0.00183571
R6356 CLK_OUT.n329 CLK_OUT.n326 0.00182678
R6357 CLK_OUT.n511 CLK_OUT.n510 0.00180952
R6358 CLK_OUT.n1223 CLK_OUT.n57 0.0017973
R6359 CLK_OUT.n1296 CLK_OUT.n1295 0.0017973
R6360 CLK_OUT.n500 CLK_OUT.n391 0.0017973
R6361 CLK_OUT.n633 CLK_OUT.n223 0.0017973
R6362 CLK_OUT.n967 CLK_OUT.n190 0.0017897
R6363 CLK_OUT.n1078 CLK_OUT.n137 0.0017897
R6364 CLK_OUT.n533 CLK_OUT.n532 0.00178256
R6365 CLK_OUT.n539 CLK_OUT.n380 0.00178256
R6366 CLK_OUT.n609 CLK_OUT.n608 0.00178256
R6367 CLK_OUT.n597 CLK_OUT.n357 0.00176044
R6368 CLK_OUT.n1162 CLK_OUT.n1161 0.00175714
R6369 CLK_OUT.n512 CLK_OUT.n389 0.00173095
R6370 CLK_OUT.n628 CLK_OUT.n627 0.00173095
R6371 CLK_OUT.n459 CLK_OUT.n458 0.00171622
R6372 CLK_OUT.n1052 CLK_OUT.n1051 0.00171347
R6373 CLK_OUT.n1190 CLK_OUT.n77 0.0016941
R6374 CLK_OUT.n1331 CLK_OUT.n1327 0.0016941
R6375 CLK_OUT.n480 CLK_OUT.n400 0.0016941
R6376 CLK_OUT.n656 CLK_OUT.n337 0.0016941
R6377 CLK_OUT.n682 CLK_OUT.n681 0.0016941
R6378 CLK_OUT.n660 CLK_OUT.n659 0.00165238
R6379 CLK_OUT.n565 CLK_OUT.n371 0.00162776
R6380 CLK_OUT.n575 CLK_OUT.n574 0.00162776
R6381 CLK_OUT.n630 CLK_OUT.n347 0.00162776
R6382 CLK_OUT.n713 CLK_OUT.n315 0.00162776
R6383 CLK_OUT.n478 CLK_OUT.n477 0.00162619
R6384 CLK_OUT.n509 CLK_OUT.n392 0.00160565
R6385 CLK_OUT.n972 CLK_OUT.n188 0.00158354
R6386 CLK_OUT.n1083 CLK_OUT.n135 0.00158354
R6387 CLK_OUT.n729 CLK_OUT.n308 0.00158354
R6388 CLK_OUT.n803 CLK_OUT.n802 0.00158354
R6389 CLK_OUT.n1251 CLK_OUT.n1250 0.00156143
R6390 CLK_OUT.n1272 CLK_OUT.n1271 0.00156143
R6391 CLK_OUT.n449 CLK_OUT.n448 0.00156143
R6392 CLK_OUT.n692 CLK_OUT.n691 0.00156143
R6393 CLK_OUT.n1054 CLK_OUT.n152 0.00156143
R6394 CLK_OUT.n1160 CLK_OUT.n101 0.00156143
R6395 CLK_OUT.n781 CLK_OUT.n780 0.00156143
R6396 CLK_OUT.n852 CLK_OUT.n274 0.00156143
R6397 CLK_OUT.n543 CLK_OUT.n542 0.00154762
R6398 CLK_OUT.n595 CLK_OUT.n594 0.00154762
R6399 CLK_OUT.n513 CLK_OUT.n390 0.00153931
R6400 CLK_OUT.n626 CLK_OUT.n349 0.00153931
R6401 CLK_OUT.n545 CLK_OUT.n544 0.00149509
R6402 CLK_OUT.n1165 CLK_OUT.n1164 0.00149509
R6403 CLK_OUT.n598 CLK_OUT.n358 0.00147297
R6404 CLK_OUT.n661 CLK_OUT.n335 0.00147297
R6405 CLK_OUT.n446 CLK_OUT.n414 0.00146905
R6406 CLK_OUT.n694 CLK_OUT.n693 0.00146905
R6407 CLK_OUT.n476 CLK_OUT.n401 0.00145086
R6408 CLK_OUT.n1209 CLK_OUT.n1208 0.00140663
R6409 CLK_OUT.n1313 CLK_OUT.n39 0.00140663
R6410 CLK_OUT.n481 CLK_OUT.n401 0.00140663
R6411 CLK_OUT.n662 CLK_OUT.n661 0.00140663
R6412 CLK_OUT.n577 CLK_OUT.n576 0.00139048
R6413 CLK_OUT.n544 CLK_OUT.n378 0.00138452
R6414 CLK_OUT.n593 CLK_OUT.n358 0.00138452
R6415 CLK_OUT.n438 CLK_OUT.n437 0.00136429
R6416 CLK_OUT.n554 CLK_OUT.n375 0.00136429
R6417 CLK_OUT.n560 CLK_OUT.n370 0.00136429
R6418 CLK_OUT.n514 CLK_OUT.n513 0.00134029
R6419 CLK_OUT.n631 CLK_OUT.n349 0.00134029
R6420 CLK_OUT.n586 CLK_OUT.n585 0.00133809
R6421 CLK_OUT.n703 CLK_OUT.n702 0.00133809
R6422 CLK_OUT.n448 CLK_OUT.n447 0.00131818
R6423 CLK_OUT.n692 CLK_OUT.n324 0.00131818
R6424 CLK_OUT.n1054 CLK_OUT.n1053 0.00131818
R6425 CLK_OUT.n743 CLK_OUT.n304 0.00129607
R6426 CLK_OUT.n765 CLK_OUT.n299 0.00129607
R6427 CLK_OUT.n820 CLK_OUT.n819 0.00129607
R6428 CLK_OUT.n843 CLK_OUT.n280 0.00129607
R6429 CLK_OUT.n461 CLK_OUT.n460 0.00128571
R6430 CLK_OUT.n679 CLK_OUT.n330 0.00128571
R6431 CLK_OUT.n1235 CLK_OUT.n56 0.00125184
R6432 CLK_OUT.n1291 CLK_OUT.n1289 0.00125184
R6433 CLK_OUT.n514 CLK_OUT.n392 0.00125184
R6434 CLK_OUT.n575 CLK_OUT.n365 0.00125184
R6435 CLK_OUT.n631 CLK_OUT.n630 0.00125184
R6436 CLK_OUT.n439 CLK_OUT.n417 0.00122973
R6437 CLK_OUT.n556 CLK_OUT.n555 0.00122973
R6438 CLK_OUT.n374 CLK_OUT.n371 0.00122973
R6439 CLK_OUT.n584 CLK_OUT.n362 0.00120762
R6440 CLK_OUT.n701 CLK_OUT.n321 0.00120762
R6441 CLK_OUT.n534 CLK_OUT.n383 0.00120714
R6442 CLK_OUT.n611 CLK_OUT.n354 0.00120714
R6443 CLK_OUT.n481 CLK_OUT.n480 0.0011855
R6444 CLK_OUT.n662 CLK_OUT.n337 0.0011855
R6445 CLK_OUT.n459 CLK_OUT.n408 0.00116339
R6446 CLK_OUT.n681 CLK_OUT.n680 0.00116339
R6447 CLK_OUT.n984 CLK_OUT.n186 0.00114865
R6448 CLK_OUT.n1095 CLK_OUT.n133 0.00114865
R6449 CLK_OUT.n733 CLK_OUT.n732 0.00114865
R6450 CLK_OUT.n807 CLK_OUT.n259 0.00114865
R6451 CLK_OUT.n651 CLK_OUT.n340 0.00112857
R6452 CLK_OUT.n598 CLK_OUT.n597 0.00111916
R6453 CLK_OUT.n494 CLK_OUT.n397 0.00110238
R6454 CLK_OUT.n1227 CLK_OUT.n1226 0.00109705
R6455 CLK_OUT.n1294 CLK_OUT.n1293 0.00109705
R6456 CLK_OUT.n533 CLK_OUT.n384 0.00109705
R6457 CLK_OUT.n545 CLK_OUT.n380 0.00109705
R6458 CLK_OUT.n610 CLK_OUT.n609 0.00109705
R6459 CLK_OUT.n1165 CLK_OUT.n100 0.00109705
R6460 CLK_OUT.n761 CLK_OUT.n760 0.00105283
R6461 CLK_OUT.n839 CLK_OUT.n838 0.00105283
R6462 CLK_OUT.n1336 CLK_OUT.n34 0.00105283
R6463 CLK_OUT.n1258 CLK_OUT.n8 0.00104054
R6464 CLK_OUT.n564 CLK_OUT.n214 0.00104054
R6465 CLK_OUT.n450 CLK_OUT.n449 0.00103071
R6466 CLK_OUT.n650 CLK_OUT.n341 0.00103071
R6467 CLK_OUT.n691 CLK_OUT.n326 0.00103071
R6468 CLK_OUT.n427 CLK_OUT.n420 0.00103071
R6469 CLK_OUT.n969 CLK_OUT.n968 0.00103071
R6470 CLK_OUT.n1080 CLK_OUT.n1079 0.00103071
R6471 CLK_OUT.n706 CLK_OUT.n319 0.00103071
R6472 CLK_OUT.n746 CLK_OUT.n745 0.00103071
R6473 CLK_OUT.n826 CLK_OUT.n825 0.00103071
R6474 CLK_OUT.n493 CLK_OUT.n492 0.0010086
R6475 CLK_OUT.n566 CLK_OUT.n565 0.000964373
R6476 CLK_OUT.n574 CLK_OUT.n367 0.000964373
R6477 CLK_OUT.n422 CLK_OUT.n421 0.000964373
R6478 CLK_OUT.n93 CLK_OUT.n90 0.000964373
R6479 CLK_OUT.n713 CLK_OUT.n316 0.000964373
R6480 CLK_OUT.n69 CLK_OUT.n66 0.00094226
R6481 CLK_OUT.n1309 CLK_OUT.n1308 0.00094226
R6482 CLK_OUT.n187 CLK_OUT.n182 0.000932432
R6483 CLK_OUT.n134 CLK_OUT.n129 0.000932432
R6484 CLK_OUT.n737 CLK_OUT.n239 0.000932432
R6485 CLK_OUT.n813 CLK_OUT.n260 0.000932432
R6486 CLK_OUT.n432 CLK_OUT.n419 0.000898034
R6487 CLK_OUT.n683 CLK_OUT.n682 0.000898034
R6488 CLK_OUT.n458 CLK_OUT.n410 0.000875921
R6489 CLK_OUT.n716 CLK_OUT.n318 0.000853808
R6490 CLK_OUT.n1152 CLK_OUT.n1151 0.000831695
R6491 CLK_OUT.n1155 CLK_OUT.n1154 0.000814286
R6492 CLK_OUT.n532 CLK_OUT.n382 0.000809582
R6493 CLK_OUT.n608 CLK_OUT.n605 0.000809582
R6494 CLK_OUT.n1244 CLK_OUT.n1243 0.000787469
R6495 CLK_OUT.n1278 CLK_OUT.n1277 0.000787469
R6496 CLK_OUT.n995 CLK_OUT.n994 0.000787469
R6497 CLK_OUT.n1106 CLK_OUT.n1105 0.000787469
R6498 CLK_OUT.n1153 CLK_OUT.n102 0.000765356
R6499 CLK_OUT.n731 CLK_OUT.n306 0.000765356
R6500 CLK_OUT.n776 CLK_OUT.n296 0.000765356
R6501 CLK_OUT.n809 CLK_OUT.n808 0.000765356
R6502 CLK_OUT.n858 CLK_OUT.n857 0.000765356
R6503 CLK_OUT.n649 CLK_OUT.n339 0.000743243
R6504 CLK_OUT.n491 CLK_OUT.n488 0.00072113
R6505 CLK_OUT.n83 CLK_OUT.n82 0.000716216
R6506 CLK_OUT.n1323 CLK_OUT.n23 0.000716216
R6507 CLK_OUT.n457 CLK_OUT.n200 0.000716216
R6508 CLK_OUT.n327 CLK_OUT.n229 0.000716216
R6509 CLK_OUT.n502 CLK_OUT.n394 0.000676904
R6510 CLK_OUT.n1194 CLK_OUT.n1193 0.000654791
R6511 CLK_OUT.n1321 CLK_OUT.n36 0.000654791
R6512 CLK_OUT.n639 CLK_OUT.n638 0.000654791
R6513 CLK_OUT.n619 CLK_OUT.n351 0.000588452
R6514 CLK_OUT.n522 CLK_OUT.n521 0.000566339
R6515 CLK_OUT.n1184 CLK_OUT.n89 0.000522113
R6516 CLK_OUT.n472 CLK_OUT.n471 0.000522113
R6517 Y0.n1376 Y0.n1373 15.1827
R6518 Y0.n1375 Y0.n1374 15.0005
R6519 Y0.n1377 Y0 10.582
R6520 Y0 Y0.n1376 9.43874
R6521 Y0.n1377 Y0 9.19322
R6522 Y0.n1369 Y0.n4 2.2505
R6523 Y0.n19 Y0.n2 2.2505
R6524 Y0.n27 Y0.n23 2.2505
R6525 Y0.n33 Y0.n26 2.2505
R6526 Y0.n1305 Y0.n29 2.2505
R6527 Y0.n1297 Y0.n1296 2.2505
R6528 Y0.n1291 Y0.n1290 2.2505
R6529 Y0.n1275 Y0.n46 2.2505
R6530 Y0.n61 Y0.n55 2.2505
R6531 Y0.n1243 Y0.n60 2.2505
R6532 Y0.n1236 Y0.n63 2.2505
R6533 Y0.n76 Y0.n72 2.2505
R6534 Y0.n1211 Y0.n74 2.2505
R6535 Y0.n94 Y0.n84 2.2505
R6536 Y0.n1192 Y0.n86 2.2505
R6537 Y0.n962 Y0.n210 2.2505
R6538 Y0.n960 Y0.n212 2.2505
R6539 Y0.n956 Y0.n215 2.2505
R6540 Y0.n954 Y0.n217 2.2505
R6541 Y0.n950 Y0.n220 2.2505
R6542 Y0.n948 Y0.n222 2.2505
R6543 Y0.n944 Y0.n225 2.2505
R6544 Y0.n942 Y0.n227 2.2505
R6545 Y0.n373 Y0.n228 2.2505
R6546 Y0.n937 Y0.n231 2.2505
R6547 Y0.n629 Y0.n233 2.2505
R6548 Y0.n931 Y0.n236 2.2505
R6549 Y0.n676 Y0.n238 2.2505
R6550 Y0.n925 Y0.n241 2.2505
R6551 Y0.n332 Y0.n243 2.2505
R6552 Y0.n963 Y0.n962 2.2505
R6553 Y0.n960 Y0.n959 2.2505
R6554 Y0.n957 Y0.n956 2.2505
R6555 Y0.n954 Y0.n953 2.2505
R6556 Y0.n951 Y0.n950 2.2505
R6557 Y0.n948 Y0.n947 2.2505
R6558 Y0.n945 Y0.n944 2.2505
R6559 Y0.n942 Y0.n941 2.2505
R6560 Y0.n940 Y0.n228 2.2505
R6561 Y0.n937 Y0.n229 2.2505
R6562 Y0.n934 Y0.n233 2.2505
R6563 Y0.n931 Y0.n234 2.2505
R6564 Y0.n928 Y0.n238 2.2505
R6565 Y0.n925 Y0.n239 2.2505
R6566 Y0.n922 Y0.n243 2.2505
R6567 Y0.n1179 Y0.n1178 2.2505
R6568 Y0.n1180 Y0.n1176 2.2505
R6569 Y0.n1175 Y0.n107 2.2505
R6570 Y0.n1174 Y0.n1173 2.2505
R6571 Y0.n109 Y0.n108 2.2505
R6572 Y0.n1132 Y0.n1131 2.2505
R6573 Y0.n1139 Y0.n1130 2.2505
R6574 Y0.n1140 Y0.n1129 2.2505
R6575 Y0.n1128 Y0.n129 2.2505
R6576 Y0.n1127 Y0.n1126 2.2505
R6577 Y0.n131 Y0.n130 2.2505
R6578 Y0.n1105 Y0.n1104 2.2505
R6579 Y0.n1103 Y0.n142 2.2505
R6580 Y0.n1102 Y0.n1101 2.2505
R6581 Y0.n144 Y0.n143 2.2505
R6582 Y0.n1078 Y0.n1077 2.2505
R6583 Y0.n1079 Y0.n1076 2.2505
R6584 Y0.n1075 Y0.n155 2.2505
R6585 Y0.n1074 Y0.n1073 2.2505
R6586 Y0.n157 Y0.n156 2.2505
R6587 Y0.n1023 Y0.n1022 2.2505
R6588 Y0.n1024 Y0.n1021 2.2505
R6589 Y0.n1025 Y0.n1020 2.2505
R6590 Y0.n1026 Y0.n1019 2.2505
R6591 Y0.n1027 Y0.n1018 2.2505
R6592 Y0.n1017 Y0.n182 2.2505
R6593 Y0.n1016 Y0.n1015 2.2505
R6594 Y0.n184 Y0.n183 2.2505
R6595 Y0.n994 Y0.n993 2.2505
R6596 Y0.n992 Y0.n195 2.2505
R6597 Y0.n991 Y0.n990 2.2505
R6598 Y0.n197 Y0.n196 2.2505
R6599 Y0.n967 Y0.n966 2.2505
R6600 Y0.n968 Y0.n965 2.2505
R6601 Y0.n969 Y0.n968 2.2505
R6602 Y0.n967 Y0.n201 2.2505
R6603 Y0.n981 Y0.n197 2.2505
R6604 Y0.n990 Y0.n989 2.2505
R6605 Y0.n199 Y0.n195 2.2505
R6606 Y0.n995 Y0.n994 2.2505
R6607 Y0.n1006 Y0.n184 2.2505
R6608 Y0.n1015 Y0.n1014 2.2505
R6609 Y0.n182 Y0.n178 2.2505
R6610 Y0.n1028 Y0.n1027 2.2505
R6611 Y0.n1026 Y0.n171 2.2505
R6612 Y0.n1025 Y0.n169 2.2505
R6613 Y0.n1024 Y0.n167 2.2505
R6614 Y0.n1023 Y0.n165 2.2505
R6615 Y0.n1054 Y0.n157 2.2505
R6616 Y0.n1073 Y0.n1072 2.2505
R6617 Y0.n1065 Y0.n155 2.2505
R6618 Y0.n1080 Y0.n1079 2.2505
R6619 Y0.n1078 Y0.n148 2.2505
R6620 Y0.n1092 Y0.n144 2.2505
R6621 Y0.n1101 Y0.n1100 2.2505
R6622 Y0.n146 Y0.n142 2.2505
R6623 Y0.n1106 Y0.n1105 2.2505
R6624 Y0.n1117 Y0.n131 2.2505
R6625 Y0.n1126 Y0.n1125 2.2505
R6626 Y0.n129 Y0.n126 2.2505
R6627 Y0.n1141 Y0.n1140 2.2505
R6628 Y0.n1139 Y0.n1138 2.2505
R6629 Y0.n1132 Y0.n117 2.2505
R6630 Y0.n1154 Y0.n109 2.2505
R6631 Y0.n1173 Y0.n1172 2.2505
R6632 Y0.n1162 Y0.n107 2.2505
R6633 Y0.n1181 Y0.n1180 2.2505
R6634 Y0.n1179 Y0.n99 2.2505
R6635 Y0.n919 Y0.n246 2.2505
R6636 Y0.n918 Y0.n247 2.2505
R6637 Y0.n917 Y0.n248 2.2505
R6638 Y0.n745 Y0.n249 2.2505
R6639 Y0.n913 Y0.n251 2.2505
R6640 Y0.n912 Y0.n252 2.2505
R6641 Y0.n911 Y0.n253 2.2505
R6642 Y0.n760 Y0.n254 2.2505
R6643 Y0.n907 Y0.n256 2.2505
R6644 Y0.n906 Y0.n257 2.2505
R6645 Y0.n905 Y0.n258 2.2505
R6646 Y0.n310 Y0.n259 2.2505
R6647 Y0.n901 Y0.n261 2.2505
R6648 Y0.n900 Y0.n262 2.2505
R6649 Y0.n899 Y0.n263 2.2505
R6650 Y0.n799 Y0.n264 2.2505
R6651 Y0.n895 Y0.n266 2.2505
R6652 Y0.n894 Y0.n267 2.2505
R6653 Y0.n893 Y0.n268 2.2505
R6654 Y0.n817 Y0.n269 2.2505
R6655 Y0.n889 Y0.n271 2.2505
R6656 Y0.n888 Y0.n272 2.2505
R6657 Y0.n887 Y0.n273 2.2505
R6658 Y0.n834 Y0.n274 2.2505
R6659 Y0.n883 Y0.n276 2.2505
R6660 Y0.n882 Y0.n277 2.2505
R6661 Y0.n881 Y0.n278 2.2505
R6662 Y0.n293 Y0.n279 2.2505
R6663 Y0.n877 Y0.n281 2.2505
R6664 Y0.n876 Y0.n282 2.2505
R6665 Y0.n875 Y0.n873 2.2505
R6666 Y0.n287 Y0.n8 2.2505
R6667 Y0.n1364 Y0.n1363 2.2505
R6668 Y0.n10 Y0.n5 2.2505
R6669 Y0.n1366 Y0.n5 2.2505
R6670 Y0.n1365 Y0.n1364 2.2505
R6671 Y0.n8 Y0.n7 2.2505
R6672 Y0.n875 Y0.n874 2.2505
R6673 Y0.n876 Y0.n280 2.2505
R6674 Y0.n878 Y0.n877 2.2505
R6675 Y0.n879 Y0.n279 2.2505
R6676 Y0.n881 Y0.n880 2.2505
R6677 Y0.n882 Y0.n275 2.2505
R6678 Y0.n884 Y0.n883 2.2505
R6679 Y0.n885 Y0.n274 2.2505
R6680 Y0.n887 Y0.n886 2.2505
R6681 Y0.n888 Y0.n270 2.2505
R6682 Y0.n890 Y0.n889 2.2505
R6683 Y0.n891 Y0.n269 2.2505
R6684 Y0.n893 Y0.n892 2.2505
R6685 Y0.n894 Y0.n265 2.2505
R6686 Y0.n896 Y0.n895 2.2505
R6687 Y0.n897 Y0.n264 2.2505
R6688 Y0.n899 Y0.n898 2.2505
R6689 Y0.n900 Y0.n260 2.2505
R6690 Y0.n902 Y0.n901 2.2505
R6691 Y0.n903 Y0.n259 2.2505
R6692 Y0.n905 Y0.n904 2.2505
R6693 Y0.n906 Y0.n255 2.2505
R6694 Y0.n908 Y0.n907 2.2505
R6695 Y0.n909 Y0.n254 2.2505
R6696 Y0.n911 Y0.n910 2.2505
R6697 Y0.n912 Y0.n250 2.2505
R6698 Y0.n914 Y0.n913 2.2505
R6699 Y0.n915 Y0.n249 2.2505
R6700 Y0.n917 Y0.n916 2.2505
R6701 Y0.n918 Y0.n245 2.2505
R6702 Y0.n920 Y0.n919 2.2505
R6703 Y0.n1369 Y0.n1 2.2505
R6704 Y0.n2 Y0.n0 2.2505
R6705 Y0.n1328 Y0.n27 2.2505
R6706 Y0.n1325 Y0.n26 2.2505
R6707 Y0.n29 Y0.n28 2.2505
R6708 Y0.n1296 Y0.n1295 2.2505
R6709 Y0.n1292 Y0.n1291 2.2505
R6710 Y0.n46 Y0.n45 2.2505
R6711 Y0.n1256 Y0.n61 2.2505
R6712 Y0.n1253 Y0.n60 2.2505
R6713 Y0.n63 Y0.n62 2.2505
R6714 Y0.n1225 Y0.n72 2.2505
R6715 Y0.n74 Y0.n73 2.2505
R6716 Y0.n1205 Y0.n84 2.2505
R6717 Y0.n86 Y0.n85 2.2505
R6718 Y0.n14 Y0.n13 2.2005
R6719 Y0.n1191 Y0.n98 2.2005
R6720 Y0.n1194 Y0.n1193 2.2005
R6721 Y0.n89 Y0.n87 2.2005
R6722 Y0.n1201 Y0.n1200 2.2005
R6723 Y0.n1199 Y0.n88 2.2005
R6724 Y0.n96 Y0.n95 2.2005
R6725 Y0.n93 Y0.n92 2.2005
R6726 Y0.n90 Y0.n83 2.2005
R6727 Y0.n1209 Y0.n80 2.2005
R6728 Y0.n1213 Y0.n1212 2.2005
R6729 Y0.n1210 Y0.n82 2.2005
R6730 Y0.n81 Y0.n75 2.2005
R6731 Y0.n1221 Y0.n1220 2.2005
R6732 Y0.n1219 Y0.n77 2.2005
R6733 Y0.n71 Y0.n70 2.2005
R6734 Y0.n1230 Y0.n1229 2.2005
R6735 Y0.n1232 Y0.n69 2.2005
R6736 Y0.n1234 Y0.n1233 2.2005
R6737 Y0.n1235 Y0.n68 2.2005
R6738 Y0.n1238 Y0.n1237 2.2005
R6739 Y0.n66 Y0.n64 2.2005
R6740 Y0.n1249 Y0.n1248 2.2005
R6741 Y0.n1247 Y0.n65 2.2005
R6742 Y0.n1245 Y0.n1244 2.2005
R6743 Y0.n59 Y0.n58 2.2005
R6744 Y0.n1262 Y0.n1261 2.2005
R6745 Y0.n1260 Y0.n56 2.2005
R6746 Y0.n1268 Y0.n1267 2.2005
R6747 Y0.n1269 Y0.n54 2.2005
R6748 Y0.n1271 Y0.n1270 2.2005
R6749 Y0.n1273 Y0.n1272 2.2005
R6750 Y0.n1274 Y0.n52 2.2005
R6751 Y0.n1277 Y0.n1276 2.2005
R6752 Y0.n49 Y0.n47 2.2005
R6753 Y0.n1289 Y0.n1288 2.2005
R6754 Y0.n50 Y0.n48 2.2005
R6755 Y0.n1282 Y0.n1281 2.2005
R6756 Y0.n1283 Y0.n42 2.2005
R6757 Y0.n1298 Y0.n41 2.2005
R6758 Y0.n1300 Y0.n1299 2.2005
R6759 Y0.n1303 Y0.n1302 2.2005
R6760 Y0.n1304 Y0.n37 2.2005
R6761 Y0.n1308 Y0.n1307 2.2005
R6762 Y0.n1306 Y0.n39 2.2005
R6763 Y0.n38 Y0.n30 2.2005
R6764 Y0.n1321 Y0.n1320 2.2005
R6765 Y0.n1319 Y0.n31 2.2005
R6766 Y0.n35 Y0.n34 2.2005
R6767 Y0.n1314 Y0.n25 2.2005
R6768 Y0.n1332 Y0.n24 2.2005
R6769 Y0.n1334 Y0.n1333 2.2005
R6770 Y0.n1336 Y0.n1335 2.2005
R6771 Y0.n1338 Y0.n1337 2.2005
R6772 Y0.n1340 Y0.n1339 2.2005
R6773 Y0.n1342 Y0.n1341 2.2005
R6774 Y0.n1345 Y0.n1344 2.2005
R6775 Y0.n1346 Y0.n18 2.2005
R6776 Y0.n1348 Y0.n1347 2.2005
R6777 Y0.n1350 Y0.n1349 2.2005
R6778 Y0.n1352 Y0.n1351 2.2005
R6779 Y0.n724 Y0.n723 2.2005
R6780 Y0.n712 Y0.n711 2.2005
R6781 Y0.n710 Y0.n709 2.2005
R6782 Y0.n703 Y0.n702 2.2005
R6783 Y0.n701 Y0.n700 2.2005
R6784 Y0.n694 Y0.n339 2.2005
R6785 Y0.n685 Y0.n343 2.2005
R6786 Y0.n687 Y0.n686 2.2005
R6787 Y0.n677 Y0.n345 2.2005
R6788 Y0.n679 Y0.n678 2.2005
R6789 Y0.n675 Y0.n674 2.2005
R6790 Y0.n667 Y0.n348 2.2005
R6791 Y0.n661 Y0.n660 2.2005
R6792 Y0.n659 Y0.n658 2.2005
R6793 Y0.n654 Y0.n653 2.2005
R6794 Y0.n652 Y0.n651 2.2005
R6795 Y0.n646 Y0.n645 2.2005
R6796 Y0.n644 Y0.n643 2.2005
R6797 Y0.n637 Y0.n360 2.2005
R6798 Y0.n631 Y0.n630 2.2005
R6799 Y0.n628 Y0.n627 2.2005
R6800 Y0.n618 Y0.n365 2.2005
R6801 Y0.n620 Y0.n619 2.2005
R6802 Y0.n613 Y0.n612 2.2005
R6803 Y0.n611 Y0.n610 2.2005
R6804 Y0.n604 Y0.n603 2.2005
R6805 Y0.n602 Y0.n601 2.2005
R6806 Y0.n595 Y0.n594 2.2005
R6807 Y0.n593 Y0.n592 2.2005
R6808 Y0.n586 Y0.n585 2.2005
R6809 Y0.n584 Y0.n583 2.2005
R6810 Y0.n577 Y0.n576 2.2005
R6811 Y0.n575 Y0.n574 2.2005
R6812 Y0.n569 Y0.n384 2.2005
R6813 Y0.n560 Y0.n388 2.2005
R6814 Y0.n562 Y0.n561 2.2005
R6815 Y0.n558 Y0.n557 2.2005
R6816 Y0.n550 Y0.n391 2.2005
R6817 Y0.n544 Y0.n543 2.2005
R6818 Y0.n542 Y0.n541 2.2005
R6819 Y0.n537 Y0.n536 2.2005
R6820 Y0.n535 Y0.n534 2.2005
R6821 Y0.n529 Y0.n528 2.2005
R6822 Y0.n527 Y0.n526 2.2005
R6823 Y0.n520 Y0.n403 2.2005
R6824 Y0.n514 Y0.n513 2.2005
R6825 Y0.n511 Y0.n510 2.2005
R6826 Y0.n501 Y0.n408 2.2005
R6827 Y0.n503 Y0.n502 2.2005
R6828 Y0.n496 Y0.n495 2.2005
R6829 Y0.n494 Y0.n493 2.2005
R6830 Y0.n487 Y0.n486 2.2005
R6831 Y0.n485 Y0.n484 2.2005
R6832 Y0.n478 Y0.n477 2.2005
R6833 Y0.n476 Y0.n475 2.2005
R6834 Y0.n470 Y0.n469 2.2005
R6835 Y0.n468 Y0.n467 2.2005
R6836 Y0.n461 Y0.n423 2.2005
R6837 Y0.n452 Y0.n427 2.2005
R6838 Y0.n454 Y0.n453 2.2005
R6839 Y0.n447 Y0.n446 2.2005
R6840 Y0.n433 Y0.n207 2.2005
R6841 Y0.n970 Y0.n206 2.2005
R6842 Y0.n972 Y0.n971 2.2005
R6843 Y0.n979 Y0.n978 2.2005
R6844 Y0.n980 Y0.n200 2.2005
R6845 Y0.n983 Y0.n982 2.2005
R6846 Y0.n985 Y0.n198 2.2005
R6847 Y0.n988 Y0.n987 2.2005
R6848 Y0.n194 Y0.n193 2.2005
R6849 Y0.n998 Y0.n996 2.2005
R6850 Y0.n189 Y0.n188 2.2005
R6851 Y0.n1005 Y0.n1004 2.2005
R6852 Y0.n1008 Y0.n1007 2.2005
R6853 Y0.n1010 Y0.n185 2.2005
R6854 Y0.n1013 Y0.n1012 2.2005
R6855 Y0.n186 Y0.n176 2.2005
R6856 Y0.n1031 Y0.n1030 2.2005
R6857 Y0.n1029 Y0.n177 2.2005
R6858 Y0.n181 Y0.n180 2.2005
R6859 Y0.n179 Y0.n172 2.2005
R6860 Y0.n1039 Y0.n1038 2.2005
R6861 Y0.n1041 Y0.n1040 2.2005
R6862 Y0.n1043 Y0.n1042 2.2005
R6863 Y0.n1045 Y0.n1044 2.2005
R6864 Y0.n1047 Y0.n1046 2.2005
R6865 Y0.n1049 Y0.n1048 2.2005
R6866 Y0.n1052 Y0.n1051 2.2005
R6867 Y0.n1053 Y0.n164 2.2005
R6868 Y0.n1057 Y0.n1055 2.2005
R6869 Y0.n160 Y0.n158 2.2005
R6870 Y0.n1071 Y0.n1070 2.2005
R6871 Y0.n1069 Y0.n159 2.2005
R6872 Y0.n1067 Y0.n1066 2.2005
R6873 Y0.n1063 Y0.n154 2.2005
R6874 Y0.n1081 Y0.n153 2.2005
R6875 Y0.n1083 Y0.n1082 2.2005
R6876 Y0.n1090 Y0.n1089 2.2005
R6877 Y0.n1091 Y0.n147 2.2005
R6878 Y0.n1094 Y0.n1093 2.2005
R6879 Y0.n1096 Y0.n145 2.2005
R6880 Y0.n1099 Y0.n1098 2.2005
R6881 Y0.n141 Y0.n140 2.2005
R6882 Y0.n1109 Y0.n1107 2.2005
R6883 Y0.n136 Y0.n135 2.2005
R6884 Y0.n1116 Y0.n1115 2.2005
R6885 Y0.n1119 Y0.n1118 2.2005
R6886 Y0.n1121 Y0.n132 2.2005
R6887 Y0.n1124 Y0.n1123 2.2005
R6888 Y0.n133 Y0.n124 2.2005
R6889 Y0.n1144 Y0.n1143 2.2005
R6890 Y0.n1142 Y0.n125 2.2005
R6891 Y0.n128 Y0.n127 2.2005
R6892 Y0.n1134 Y0.n1133 2.2005
R6893 Y0.n1137 Y0.n1136 2.2005
R6894 Y0.n1135 Y0.n118 2.2005
R6895 Y0.n1152 Y0.n1151 2.2005
R6896 Y0.n1153 Y0.n116 2.2005
R6897 Y0.n1156 Y0.n1155 2.2005
R6898 Y0.n114 Y0.n110 2.2005
R6899 Y0.n1171 Y0.n1170 2.2005
R6900 Y0.n113 Y0.n111 2.2005
R6901 Y0.n1164 Y0.n1163 2.2005
R6902 Y0.n106 Y0.n104 2.2005
R6903 Y0.n1184 Y0.n1183 2.2005
R6904 Y0.n1182 Y0.n105 2.2005
R6905 Y0.n726 Y0.n725 2.2005
R6906 Y0.n735 Y0.n734 2.2005
R6907 Y0.n737 Y0.n736 2.2005
R6908 Y0.n739 Y0.n738 2.2005
R6909 Y0.n741 Y0.n740 2.2005
R6910 Y0.n742 Y0.n319 2.2005
R6911 Y0.n744 Y0.n743 2.2005
R6912 Y0.n747 Y0.n746 2.2005
R6913 Y0.n749 Y0.n748 2.2005
R6914 Y0.n751 Y0.n750 2.2005
R6915 Y0.n753 Y0.n752 2.2005
R6916 Y0.n755 Y0.n754 2.2005
R6917 Y0.n756 Y0.n315 2.2005
R6918 Y0.n759 Y0.n758 2.2005
R6919 Y0.n761 Y0.n314 2.2005
R6920 Y0.n763 Y0.n762 2.2005
R6921 Y0.n766 Y0.n765 2.2005
R6922 Y0.n764 Y0.n312 2.2005
R6923 Y0.n774 Y0.n773 2.2005
R6924 Y0.n776 Y0.n775 2.2005
R6925 Y0.n778 Y0.n777 2.2005
R6926 Y0.n780 Y0.n779 2.2005
R6927 Y0.n782 Y0.n781 2.2005
R6928 Y0.n784 Y0.n783 2.2005
R6929 Y0.n786 Y0.n785 2.2005
R6930 Y0.n788 Y0.n787 2.2005
R6931 Y0.n790 Y0.n789 2.2005
R6932 Y0.n792 Y0.n791 2.2005
R6933 Y0.n306 Y0.n305 2.2005
R6934 Y0.n798 Y0.n797 2.2005
R6935 Y0.n800 Y0.n304 2.2005
R6936 Y0.n802 Y0.n801 2.2005
R6937 Y0.n804 Y0.n803 2.2005
R6938 Y0.n806 Y0.n805 2.2005
R6939 Y0.n808 Y0.n807 2.2005
R6940 Y0.n810 Y0.n809 2.2005
R6941 Y0.n302 Y0.n301 2.2005
R6942 Y0.n816 Y0.n815 2.2005
R6943 Y0.n818 Y0.n300 2.2005
R6944 Y0.n820 Y0.n819 2.2005
R6945 Y0.n823 Y0.n822 2.2005
R6946 Y0.n825 Y0.n824 2.2005
R6947 Y0.n827 Y0.n826 2.2005
R6948 Y0.n298 Y0.n297 2.2005
R6949 Y0.n833 Y0.n832 2.2005
R6950 Y0.n835 Y0.n296 2.2005
R6951 Y0.n837 Y0.n836 2.2005
R6952 Y0.n840 Y0.n839 2.2005
R6953 Y0.n842 Y0.n841 2.2005
R6954 Y0.n845 Y0.n844 2.2005
R6955 Y0.n843 Y0.n294 2.2005
R6956 Y0.n852 Y0.n851 2.2005
R6957 Y0.n854 Y0.n853 2.2005
R6958 Y0.n856 Y0.n855 2.2005
R6959 Y0.n858 Y0.n857 2.2005
R6960 Y0.n860 Y0.n859 2.2005
R6961 Y0.n862 Y0.n861 2.2005
R6962 Y0.n864 Y0.n863 2.2005
R6963 Y0.n285 Y0.n283 2.2005
R6964 Y0.n872 Y0.n871 2.2005
R6965 Y0.n870 Y0.n284 2.2005
R6966 Y0.n289 Y0.n288 2.2005
R6967 Y0.n286 Y0.n9 2.2005
R6968 Y0.n1362 Y0.n1361 2.2005
R6969 Y0.n1360 Y0.n11 2.2005
R6970 Y0.n1370 Y0.n3 1.8005
R6971 Y0.n1326 Y0.n21 1.8005
R6972 Y0.n1331 Y0.n1330 1.8005
R6973 Y0.n1323 Y0.n1322 1.8005
R6974 Y0.n44 Y0.n40 1.8005
R6975 Y0.n1280 Y0.n43 1.8005
R6976 Y0.n1254 Y0.n53 1.8005
R6977 Y0.n1259 Y0.n1258 1.8005
R6978 Y0.n1251 Y0.n1250 1.8005
R6979 Y0.n1228 Y0.n1227 1.8005
R6980 Y0.n1223 Y0.n1222 1.8005
R6981 Y0.n1208 Y0.n1207 1.8005
R6982 Y0.n1203 Y0.n1202 1.8005
R6983 Y0.n961 Y0.n211 1.8005
R6984 Y0.n416 Y0.n213 1.8005
R6985 Y0.n955 Y0.n216 1.8005
R6986 Y0.n512 Y0.n218 1.8005
R6987 Y0.n949 Y0.n221 1.8005
R6988 Y0.n559 Y0.n223 1.8005
R6989 Y0.n943 Y0.n226 1.8005
R6990 Y0.n938 Y0.n230 1.8005
R6991 Y0.n936 Y0.n232 1.8005
R6992 Y0.n932 Y0.n235 1.8005
R6993 Y0.n930 Y0.n237 1.8005
R6994 Y0.n926 Y0.n240 1.8005
R6995 Y0.n924 Y0.n242 1.8005
R6996 Y0.n961 Y0.n209 1.8005
R6997 Y0.n958 Y0.n213 1.8005
R6998 Y0.n955 Y0.n214 1.8005
R6999 Y0.n952 Y0.n218 1.8005
R7000 Y0.n949 Y0.n219 1.8005
R7001 Y0.n946 Y0.n223 1.8005
R7002 Y0.n943 Y0.n224 1.8005
R7003 Y0.n939 Y0.n938 1.8005
R7004 Y0.n936 Y0.n935 1.8005
R7005 Y0.n933 Y0.n932 1.8005
R7006 Y0.n930 Y0.n929 1.8005
R7007 Y0.n927 Y0.n926 1.8005
R7008 Y0.n924 Y0.n923 1.8005
R7009 Y0.n1177 Y0.n100 1.8005
R7010 Y0.n1190 Y0.n100 1.8005
R7011 Y0.n1368 Y0.n6 1.8005
R7012 Y0.n1368 Y0.n1367 1.8005
R7013 Y0.n1371 Y0.n1370 1.8005
R7014 Y0.n1327 Y0.n1326 1.8005
R7015 Y0.n1330 Y0.n1329 1.8005
R7016 Y0.n1324 Y0.n1323 1.8005
R7017 Y0.n1294 Y0.n44 1.8005
R7018 Y0.n1293 Y0.n43 1.8005
R7019 Y0.n1255 Y0.n1254 1.8005
R7020 Y0.n1258 Y0.n1257 1.8005
R7021 Y0.n1252 Y0.n1251 1.8005
R7022 Y0.n1227 Y0.n1226 1.8005
R7023 Y0.n1224 Y0.n1223 1.8005
R7024 Y0.n1207 Y0.n1206 1.8005
R7025 Y0.n1204 Y0.n1203 1.8005
R7026 Y0.n964 Y0.n208 1.5005
R7027 Y0.n445 Y0.n208 1.5005
R7028 Y0.n727 Y0.n244 1.5005
R7029 Y0.n921 Y0.n244 1.5005
R7030 Y0.n731 Y0.n327 1.1125
R7031 Y0.n1169 Y0.n1168 1.10836
R7032 Y0.n1161 Y0.n112 1.10443
R7033 Y0.n1187 Y0.n102 1.10381
R7034 Y0.n730 Y0.n328 1.10372
R7035 Y0.n1157 Y0.n115 1.10339
R7036 Y0.n1164 Y0.n103 1.10272
R7037 Y0.n1167 Y0.n113 1.10272
R7038 Y0.n1160 Y0.n114 1.10272
R7039 Y0.n734 Y0.n733 1.10263
R7040 Y0.n737 Y0.n326 1.10263
R7041 Y0.n1354 Y0.n1353 1.1005
R7042 Y0.n1196 Y0.n1195 1.1005
R7043 Y0.n1198 Y0.n1197 1.1005
R7044 Y0.n91 Y0.n79 1.1005
R7045 Y0.n1215 Y0.n1214 1.1005
R7046 Y0.n1216 Y0.n78 1.1005
R7047 Y0.n1218 Y0.n1217 1.1005
R7048 Y0.n1231 Y0.n67 1.1005
R7049 Y0.n1240 Y0.n1239 1.1005
R7050 Y0.n1242 Y0.n1241 1.1005
R7051 Y0.n1246 Y0.n57 1.1005
R7052 Y0.n1264 Y0.n1263 1.1005
R7053 Y0.n1266 Y0.n1265 1.1005
R7054 Y0.n1272 Y0.n51 1.1005
R7055 Y0.n1279 Y0.n1278 1.1005
R7056 Y0.n1287 Y0.n1286 1.1005
R7057 Y0.n1285 Y0.n1284 1.1005
R7058 Y0.n1301 Y0.n36 1.1005
R7059 Y0.n1310 Y0.n1309 1.1005
R7060 Y0.n1311 Y0.n32 1.1005
R7061 Y0.n1318 Y0.n1317 1.1005
R7062 Y0.n1316 Y0.n1315 1.1005
R7063 Y0.n1313 Y0.n22 1.1005
R7064 Y0.n1312 Y0.n20 1.1005
R7065 Y0.n1343 Y0.n17 1.1005
R7066 Y0.n101 Y0.n97 1.1005
R7067 Y0.n973 Y0.n204 1.1005
R7068 Y0.n999 Y0.n191 1.1005
R7069 Y0.n1058 Y0.n162 1.1005
R7070 Y0.n1084 Y0.n151 1.1005
R7071 Y0.n1110 Y0.n138 1.1005
R7072 Y0.n1186 Y0.n1185 1.1005
R7073 Y0.n1166 Y0.n1165 1.1005
R7074 Y0.n1159 Y0.n1158 1.1005
R7075 Y0.n1150 Y0.n1149 1.1005
R7076 Y0.n1146 Y0.n1145 1.1005
R7077 Y0.n1112 Y0.n1111 1.1005
R7078 Y0.n1088 Y0.n1087 1.1005
R7079 Y0.n1086 Y0.n1085 1.1005
R7080 Y0.n1062 Y0.n1061 1.1005
R7081 Y0.n1060 Y0.n1059 1.1005
R7082 Y0.n1035 Y0.n168 1.1005
R7083 Y0.n1033 Y0.n1032 1.1005
R7084 Y0.n1001 Y0.n1000 1.1005
R7085 Y0.n977 Y0.n976 1.1005
R7086 Y0.n975 Y0.n974 1.1005
R7087 Y0.n442 Y0.n435 1.1005
R7088 Y0.n441 Y0.n432 1.1005
R7089 Y0.n434 Y0.n205 1.1005
R7090 Y0.n444 Y0.n443 1.1005
R7091 Y0.n723 Y0.n722 1.1005
R7092 Y0.n714 Y0.n713 1.1005
R7093 Y0.n712 Y0.n334 1.1005
R7094 Y0.n709 Y0.n708 1.1005
R7095 Y0.n705 Y0.n704 1.1005
R7096 Y0.n698 Y0.n341 1.1005
R7097 Y0.n700 Y0.n699 1.1005
R7098 Y0.n697 Y0.n340 1.1005
R7099 Y0.n692 Y0.n691 1.1005
R7100 Y0.n681 Y0.n680 1.1005
R7101 Y0.n679 Y0.n346 1.1005
R7102 Y0.n671 Y0.n347 1.1005
R7103 Y0.n669 Y0.n668 1.1005
R7104 Y0.n667 Y0.n350 1.1005
R7105 Y0.n666 Y0.n665 1.1005
R7106 Y0.n353 Y0.n352 1.1005
R7107 Y0.n648 Y0.n357 1.1005
R7108 Y0.n647 Y0.n646 1.1005
R7109 Y0.n359 Y0.n358 1.1005
R7110 Y0.n639 Y0.n638 1.1005
R7111 Y0.n637 Y0.n362 1.1005
R7112 Y0.n636 Y0.n635 1.1005
R7113 Y0.n633 Y0.n632 1.1005
R7114 Y0.n627 Y0.n364 1.1005
R7115 Y0.n624 Y0.n365 1.1005
R7116 Y0.n621 Y0.n366 1.1005
R7117 Y0.n615 Y0.n367 1.1005
R7118 Y0.n614 Y0.n613 1.1005
R7119 Y0.n369 Y0.n368 1.1005
R7120 Y0.n606 Y0.n605 1.1005
R7121 Y0.n597 Y0.n596 1.1005
R7122 Y0.n595 Y0.n375 1.1005
R7123 Y0.n592 Y0.n591 1.1005
R7124 Y0.n588 Y0.n587 1.1005
R7125 Y0.n581 Y0.n381 1.1005
R7126 Y0.n583 Y0.n582 1.1005
R7127 Y0.n580 Y0.n380 1.1005
R7128 Y0.n572 Y0.n386 1.1005
R7129 Y0.n567 Y0.n566 1.1005
R7130 Y0.n565 Y0.n388 1.1005
R7131 Y0.n562 Y0.n389 1.1005
R7132 Y0.n556 Y0.n555 1.1005
R7133 Y0.n552 Y0.n551 1.1005
R7134 Y0.n550 Y0.n393 1.1005
R7135 Y0.n549 Y0.n548 1.1005
R7136 Y0.n396 Y0.n395 1.1005
R7137 Y0.n531 Y0.n400 1.1005
R7138 Y0.n530 Y0.n529 1.1005
R7139 Y0.n402 Y0.n401 1.1005
R7140 Y0.n522 Y0.n521 1.1005
R7141 Y0.n520 Y0.n405 1.1005
R7142 Y0.n519 Y0.n518 1.1005
R7143 Y0.n516 Y0.n515 1.1005
R7144 Y0.n510 Y0.n407 1.1005
R7145 Y0.n507 Y0.n408 1.1005
R7146 Y0.n504 Y0.n409 1.1005
R7147 Y0.n498 Y0.n410 1.1005
R7148 Y0.n497 Y0.n496 1.1005
R7149 Y0.n412 Y0.n411 1.1005
R7150 Y0.n489 Y0.n488 1.1005
R7151 Y0.n487 Y0.n414 1.1005
R7152 Y0.n481 Y0.n415 1.1005
R7153 Y0.n480 Y0.n417 1.1005
R7154 Y0.n479 Y0.n478 1.1005
R7155 Y0.n475 Y0.n474 1.1005
R7156 Y0.n472 Y0.n471 1.1005
R7157 Y0.n465 Y0.n425 1.1005
R7158 Y0.n467 Y0.n466 1.1005
R7159 Y0.n464 Y0.n424 1.1005
R7160 Y0.n459 Y0.n458 1.1005
R7161 Y0.n449 Y0.n429 1.1005
R7162 Y0.n448 Y0.n447 1.1005
R7163 Y0.n439 Y0.n438 1.1005
R7164 Y0.n440 Y0.n439 1.1005
R7165 Y0.n437 Y0.n432 1.1005
R7166 Y0.n431 Y0.n430 1.1005
R7167 Y0.n457 Y0.n427 1.1005
R7168 Y0.n456 Y0.n455 1.1005
R7169 Y0.n454 Y0.n428 1.1005
R7170 Y0.n451 Y0.n450 1.1005
R7171 Y0.n460 Y0.n426 1.1005
R7172 Y0.n463 Y0.n462 1.1005
R7173 Y0.n422 Y0.n421 1.1005
R7174 Y0.n473 Y0.n420 1.1005
R7175 Y0.n419 Y0.n418 1.1005
R7176 Y0.n483 Y0.n482 1.1005
R7177 Y0.n490 Y0.n413 1.1005
R7178 Y0.n492 Y0.n491 1.1005
R7179 Y0.n500 Y0.n499 1.1005
R7180 Y0.n506 Y0.n505 1.1005
R7181 Y0.n509 Y0.n508 1.1005
R7182 Y0.n517 Y0.n406 1.1005
R7183 Y0.n523 Y0.n404 1.1005
R7184 Y0.n525 Y0.n524 1.1005
R7185 Y0.n533 Y0.n532 1.1005
R7186 Y0.n541 Y0.n540 1.1005
R7187 Y0.n539 Y0.n397 1.1005
R7188 Y0.n538 Y0.n537 1.1005
R7189 Y0.n399 Y0.n398 1.1005
R7190 Y0.n546 Y0.n545 1.1005
R7191 Y0.n547 Y0.n394 1.1005
R7192 Y0.n553 Y0.n392 1.1005
R7193 Y0.n554 Y0.n390 1.1005
R7194 Y0.n564 Y0.n563 1.1005
R7195 Y0.n574 Y0.n573 1.1005
R7196 Y0.n571 Y0.n385 1.1005
R7197 Y0.n570 Y0.n569 1.1005
R7198 Y0.n568 Y0.n387 1.1005
R7199 Y0.n383 Y0.n382 1.1005
R7200 Y0.n579 Y0.n578 1.1005
R7201 Y0.n379 Y0.n378 1.1005
R7202 Y0.n589 Y0.n377 1.1005
R7203 Y0.n590 Y0.n376 1.1005
R7204 Y0.n604 Y0.n371 1.1005
R7205 Y0.n599 Y0.n372 1.1005
R7206 Y0.n601 Y0.n600 1.1005
R7207 Y0.n598 Y0.n374 1.1005
R7208 Y0.n607 Y0.n370 1.1005
R7209 Y0.n609 Y0.n608 1.1005
R7210 Y0.n617 Y0.n616 1.1005
R7211 Y0.n623 Y0.n622 1.1005
R7212 Y0.n626 Y0.n625 1.1005
R7213 Y0.n634 Y0.n363 1.1005
R7214 Y0.n640 Y0.n361 1.1005
R7215 Y0.n642 Y0.n641 1.1005
R7216 Y0.n650 Y0.n649 1.1005
R7217 Y0.n658 Y0.n657 1.1005
R7218 Y0.n656 Y0.n354 1.1005
R7219 Y0.n655 Y0.n654 1.1005
R7220 Y0.n356 Y0.n355 1.1005
R7221 Y0.n663 Y0.n662 1.1005
R7222 Y0.n664 Y0.n351 1.1005
R7223 Y0.n670 Y0.n349 1.1005
R7224 Y0.n673 Y0.n672 1.1005
R7225 Y0.n682 Y0.n345 1.1005
R7226 Y0.n690 Y0.n343 1.1005
R7227 Y0.n689 Y0.n688 1.1005
R7228 Y0.n687 Y0.n344 1.1005
R7229 Y0.n684 Y0.n683 1.1005
R7230 Y0.n693 Y0.n342 1.1005
R7231 Y0.n696 Y0.n695 1.1005
R7232 Y0.n338 Y0.n337 1.1005
R7233 Y0.n706 Y0.n336 1.1005
R7234 Y0.n707 Y0.n335 1.1005
R7235 Y0.n715 Y0.n333 1.1005
R7236 Y0.n721 Y0.n330 1.1005
R7237 Y0.n331 Y0.n329 1.1005
R7238 Y0.n718 Y0.n717 1.1005
R7239 Y0.n1358 Y0.n1357 1.1005
R7240 Y0.n1356 Y0.n16 1.1005
R7241 Y0.n1355 Y0.n16 1.1005
R7242 Y0.n720 Y0.n331 1.1005
R7243 Y0.n719 Y0.n718 1.1005
R7244 Y0.n1359 Y0.n15 1.1005
R7245 Y0.n867 Y0.n12 1.1005
R7246 Y0.n869 Y0.n868 1.1005
R7247 Y0.n866 Y0.n865 1.1005
R7248 Y0.n291 Y0.n290 1.1005
R7249 Y0.n848 Y0.n292 1.1005
R7250 Y0.n850 Y0.n849 1.1005
R7251 Y0.n847 Y0.n846 1.1005
R7252 Y0.n838 Y0.n295 1.1005
R7253 Y0.n831 Y0.n830 1.1005
R7254 Y0.n829 Y0.n828 1.1005
R7255 Y0.n821 Y0.n299 1.1005
R7256 Y0.n814 Y0.n813 1.1005
R7257 Y0.n812 Y0.n811 1.1005
R7258 Y0.n803 Y0.n303 1.1005
R7259 Y0.n796 Y0.n795 1.1005
R7260 Y0.n794 Y0.n793 1.1005
R7261 Y0.n308 Y0.n307 1.1005
R7262 Y0.n769 Y0.n309 1.1005
R7263 Y0.n770 Y0.n311 1.1005
R7264 Y0.n772 Y0.n771 1.1005
R7265 Y0.n768 Y0.n767 1.1005
R7266 Y0.n757 Y0.n313 1.1005
R7267 Y0.n322 Y0.n316 1.1005
R7268 Y0.n323 Y0.n317 1.1005
R7269 Y0.n324 Y0.n318 1.1005
R7270 Y0.n325 Y0.n320 1.1005
R7271 Y0.n732 Y0.n321 1.1005
R7272 Y0.n729 Y0.n728 1.1005
R7273 Y0.n445 Y0.n444 0.733833
R7274 Y0.n1190 Y0.n1189 0.733833
R7275 Y0.n1359 Y0.n6 0.733833
R7276 Y0.n728 Y0.n727 0.733833
R7277 Y0.n1108 Y0.n138 0.573769
R7278 Y0.n997 Y0.n191 0.573769
R7279 Y0.n151 Y0.n149 0.573695
R7280 Y0.n204 Y0.n202 0.573695
R7281 Y0.n1056 Y0.n162 0.573346
R7282 Y0.n436 Y0.n432 0.550549
R7283 Y0.n716 Y0.n331 0.550549
R7284 Y0 Y0.n1372 0.45425
R7285 Y0.n1112 Y0.n137 0.39244
R7286 Y0.n1001 Y0.n190 0.39244
R7287 Y0.n1086 Y0.n150 0.389994
R7288 Y0.n975 Y0.n203 0.389994
R7289 Y0.n1060 Y0.n161 0.387191
R7290 Y0.n1148 Y0.n119 0.384705
R7291 Y0.n1037 Y0.n1036 0.384705
R7292 Y0.n1113 Y0.n134 0.384705
R7293 Y0.n1002 Y0.n187 0.384705
R7294 Y0.n1147 Y0.n122 0.382331
R7295 Y0.n1034 Y0.n174 0.382331
R7296 Y0.n1120 Y0.n123 0.382034
R7297 Y0.n1009 Y0.n175 0.382034
R7298 Y0.n1095 Y0.n139 0.379547
R7299 Y0.n1050 Y0.n163 0.379547
R7300 Y0.n984 Y0.n192 0.379547
R7301 Y0.n1064 Y0.n152 0.376968
R7302 Y0.n1068 Y0.n152 0.376876
R7303 Y0.n1097 Y0.n139 0.375976
R7304 Y0.n986 Y0.n192 0.375976
R7305 Y0.n166 Y0.n163 0.375884
R7306 Y0.n1122 Y0.n123 0.374982
R7307 Y0.n1011 Y0.n175 0.374982
R7308 Y0.n1147 Y0.n121 0.374889
R7309 Y0.n1034 Y0.n173 0.374889
R7310 Y0.n1148 Y0.n120 0.373984
R7311 Y0.n1036 Y0.n170 0.373984
R7312 Y0.n1114 Y0.n1113 0.373891
R7313 Y0.n1003 Y0.n1002 0.373891
R7314 Y0.n1189 Y0.n1188 0.275034
R7315 Y0.n1376 Y0.n1375 0.189306
R7316 Y0.n1375 Y0 0.0513955
R7317 Y0.n1203 Y0.n86 0.0405
R7318 Y0.n1203 Y0.n84 0.0405
R7319 Y0.n1207 Y0.n84 0.0405
R7320 Y0.n1207 Y0.n74 0.0405
R7321 Y0.n1223 Y0.n74 0.0405
R7322 Y0.n1223 Y0.n72 0.0405
R7323 Y0.n1227 Y0.n72 0.0405
R7324 Y0.n1227 Y0.n63 0.0405
R7325 Y0.n1251 Y0.n63 0.0405
R7326 Y0.n1251 Y0.n60 0.0405
R7327 Y0.n1258 Y0.n60 0.0405
R7328 Y0.n1258 Y0.n61 0.0405
R7329 Y0.n1254 Y0.n61 0.0405
R7330 Y0.n1254 Y0.n46 0.0405
R7331 Y0.n1291 Y0.n43 0.0405
R7332 Y0.n1296 Y0.n43 0.0405
R7333 Y0.n1296 Y0.n44 0.0405
R7334 Y0.n44 Y0.n29 0.0405
R7335 Y0.n1323 Y0.n29 0.0405
R7336 Y0.n1323 Y0.n26 0.0405
R7337 Y0.n1330 Y0.n26 0.0405
R7338 Y0.n1330 Y0.n27 0.0405
R7339 Y0.n1326 Y0.n27 0.0405
R7340 Y0.n1326 Y0.n2 0.0405
R7341 Y0.n1370 Y0.n2 0.0405
R7342 Y0.n1370 Y0.n1369 0.0405
R7343 Y0.n962 Y0.n961 0.0405
R7344 Y0.n961 Y0.n960 0.0405
R7345 Y0.n960 Y0.n213 0.0405
R7346 Y0.n956 Y0.n213 0.0405
R7347 Y0.n956 Y0.n955 0.0405
R7348 Y0.n955 Y0.n954 0.0405
R7349 Y0.n954 Y0.n218 0.0405
R7350 Y0.n950 Y0.n218 0.0405
R7351 Y0.n950 Y0.n949 0.0405
R7352 Y0.n949 Y0.n948 0.0405
R7353 Y0.n948 Y0.n223 0.0405
R7354 Y0.n944 Y0.n223 0.0405
R7355 Y0.n944 Y0.n943 0.0405
R7356 Y0.n943 Y0.n942 0.0405
R7357 Y0.n938 Y0.n228 0.0405
R7358 Y0.n938 Y0.n937 0.0405
R7359 Y0.n937 Y0.n936 0.0405
R7360 Y0.n936 Y0.n233 0.0405
R7361 Y0.n932 Y0.n233 0.0405
R7362 Y0.n932 Y0.n931 0.0405
R7363 Y0.n931 Y0.n930 0.0405
R7364 Y0.n930 Y0.n238 0.0405
R7365 Y0.n926 Y0.n238 0.0405
R7366 Y0.n926 Y0.n925 0.0405
R7367 Y0.n925 Y0.n924 0.0405
R7368 Y0.n924 Y0.n243 0.0405
R7369 Y0.n963 Y0.n209 0.0405
R7370 Y0.n959 Y0.n209 0.0405
R7371 Y0.n959 Y0.n958 0.0405
R7372 Y0.n958 Y0.n957 0.0405
R7373 Y0.n957 Y0.n214 0.0405
R7374 Y0.n953 Y0.n214 0.0405
R7375 Y0.n953 Y0.n952 0.0405
R7376 Y0.n952 Y0.n951 0.0405
R7377 Y0.n951 Y0.n219 0.0405
R7378 Y0.n947 Y0.n219 0.0405
R7379 Y0.n947 Y0.n946 0.0405
R7380 Y0.n946 Y0.n945 0.0405
R7381 Y0.n945 Y0.n224 0.0405
R7382 Y0.n941 Y0.n224 0.0405
R7383 Y0.n940 Y0.n939 0.0405
R7384 Y0.n939 Y0.n229 0.0405
R7385 Y0.n935 Y0.n229 0.0405
R7386 Y0.n935 Y0.n934 0.0405
R7387 Y0.n934 Y0.n933 0.0405
R7388 Y0.n933 Y0.n234 0.0405
R7389 Y0.n929 Y0.n234 0.0405
R7390 Y0.n929 Y0.n928 0.0405
R7391 Y0.n928 Y0.n927 0.0405
R7392 Y0.n927 Y0.n239 0.0405
R7393 Y0.n923 Y0.n239 0.0405
R7394 Y0.n923 Y0.n922 0.0405
R7395 Y0.n1204 Y0.n85 0.0405
R7396 Y0.n1205 Y0.n1204 0.0405
R7397 Y0.n1206 Y0.n1205 0.0405
R7398 Y0.n1206 Y0.n73 0.0405
R7399 Y0.n1224 Y0.n73 0.0405
R7400 Y0.n1225 Y0.n1224 0.0405
R7401 Y0.n1226 Y0.n1225 0.0405
R7402 Y0.n1226 Y0.n62 0.0405
R7403 Y0.n1252 Y0.n62 0.0405
R7404 Y0.n1253 Y0.n1252 0.0405
R7405 Y0.n1257 Y0.n1253 0.0405
R7406 Y0.n1257 Y0.n1256 0.0405
R7407 Y0.n1256 Y0.n1255 0.0405
R7408 Y0.n1255 Y0.n45 0.0405
R7409 Y0.n1293 Y0.n1292 0.0405
R7410 Y0.n1295 Y0.n1293 0.0405
R7411 Y0.n1295 Y0.n1294 0.0405
R7412 Y0.n1294 Y0.n28 0.0405
R7413 Y0.n1324 Y0.n28 0.0405
R7414 Y0.n1325 Y0.n1324 0.0405
R7415 Y0.n1329 Y0.n1325 0.0405
R7416 Y0.n1329 Y0.n1328 0.0405
R7417 Y0.n1328 Y0.n1327 0.0405
R7418 Y0.n1327 Y0.n0 0.0405
R7419 Y0.n1371 Y0.n1 0.0405
R7420 Y0.n1372 Y0.n1371 0.0386622
R7421 Y0.n1291 Y0.n46 0.0360676
R7422 Y0.n942 Y0.n228 0.0360676
R7423 Y0.n941 Y0.n940 0.0360676
R7424 Y0.n966 Y0.n965 0.0360676
R7425 Y0.n966 Y0.n196 0.0360676
R7426 Y0.n991 Y0.n196 0.0360676
R7427 Y0.n992 Y0.n991 0.0360676
R7428 Y0.n993 Y0.n992 0.0360676
R7429 Y0.n993 Y0.n183 0.0360676
R7430 Y0.n1016 Y0.n183 0.0360676
R7431 Y0.n1017 Y0.n1016 0.0360676
R7432 Y0.n1018 Y0.n1017 0.0360676
R7433 Y0.n1019 Y0.n1018 0.0360676
R7434 Y0.n1020 Y0.n1019 0.0360676
R7435 Y0.n1021 Y0.n1020 0.0360676
R7436 Y0.n1022 Y0.n1021 0.0360676
R7437 Y0.n1022 Y0.n156 0.0360676
R7438 Y0.n1074 Y0.n156 0.0360676
R7439 Y0.n1075 Y0.n1074 0.0360676
R7440 Y0.n1076 Y0.n1075 0.0360676
R7441 Y0.n1077 Y0.n1076 0.0360676
R7442 Y0.n1077 Y0.n143 0.0360676
R7443 Y0.n1102 Y0.n143 0.0360676
R7444 Y0.n1103 Y0.n1102 0.0360676
R7445 Y0.n1104 Y0.n1103 0.0360676
R7446 Y0.n1104 Y0.n130 0.0360676
R7447 Y0.n1127 Y0.n130 0.0360676
R7448 Y0.n1128 Y0.n1127 0.0360676
R7449 Y0.n1129 Y0.n1128 0.0360676
R7450 Y0.n1130 Y0.n1129 0.0360676
R7451 Y0.n1131 Y0.n1130 0.0360676
R7452 Y0.n1131 Y0.n108 0.0360676
R7453 Y0.n1174 Y0.n108 0.0360676
R7454 Y0.n1175 Y0.n1174 0.0360676
R7455 Y0.n1176 Y0.n1175 0.0360676
R7456 Y0.n1178 Y0.n1176 0.0360676
R7457 Y0.n968 Y0.n967 0.0360676
R7458 Y0.n967 Y0.n197 0.0360676
R7459 Y0.n990 Y0.n197 0.0360676
R7460 Y0.n990 Y0.n195 0.0360676
R7461 Y0.n994 Y0.n195 0.0360676
R7462 Y0.n994 Y0.n184 0.0360676
R7463 Y0.n1015 Y0.n184 0.0360676
R7464 Y0.n1015 Y0.n182 0.0360676
R7465 Y0.n1027 Y0.n182 0.0360676
R7466 Y0.n1027 Y0.n1026 0.0360676
R7467 Y0.n1026 Y0.n1025 0.0360676
R7468 Y0.n1025 Y0.n1024 0.0360676
R7469 Y0.n1024 Y0.n1023 0.0360676
R7470 Y0.n1023 Y0.n157 0.0360676
R7471 Y0.n1073 Y0.n157 0.0360676
R7472 Y0.n1073 Y0.n155 0.0360676
R7473 Y0.n1079 Y0.n155 0.0360676
R7474 Y0.n1079 Y0.n1078 0.0360676
R7475 Y0.n1078 Y0.n144 0.0360676
R7476 Y0.n1101 Y0.n144 0.0360676
R7477 Y0.n1101 Y0.n142 0.0360676
R7478 Y0.n1105 Y0.n142 0.0360676
R7479 Y0.n1105 Y0.n131 0.0360676
R7480 Y0.n1126 Y0.n131 0.0360676
R7481 Y0.n1126 Y0.n129 0.0360676
R7482 Y0.n1140 Y0.n129 0.0360676
R7483 Y0.n1140 Y0.n1139 0.0360676
R7484 Y0.n1139 Y0.n1132 0.0360676
R7485 Y0.n1132 Y0.n109 0.0360676
R7486 Y0.n1173 Y0.n109 0.0360676
R7487 Y0.n1173 Y0.n107 0.0360676
R7488 Y0.n1180 Y0.n107 0.0360676
R7489 Y0.n1180 Y0.n1179 0.0360676
R7490 Y0.n919 Y0.n918 0.0360676
R7491 Y0.n918 Y0.n917 0.0360676
R7492 Y0.n917 Y0.n249 0.0360676
R7493 Y0.n913 Y0.n249 0.0360676
R7494 Y0.n913 Y0.n912 0.0360676
R7495 Y0.n912 Y0.n911 0.0360676
R7496 Y0.n911 Y0.n254 0.0360676
R7497 Y0.n907 Y0.n254 0.0360676
R7498 Y0.n907 Y0.n906 0.0360676
R7499 Y0.n906 Y0.n905 0.0360676
R7500 Y0.n905 Y0.n259 0.0360676
R7501 Y0.n901 Y0.n259 0.0360676
R7502 Y0.n901 Y0.n900 0.0360676
R7503 Y0.n900 Y0.n899 0.0360676
R7504 Y0.n899 Y0.n264 0.0360676
R7505 Y0.n895 Y0.n264 0.0360676
R7506 Y0.n895 Y0.n894 0.0360676
R7507 Y0.n894 Y0.n893 0.0360676
R7508 Y0.n893 Y0.n269 0.0360676
R7509 Y0.n889 Y0.n269 0.0360676
R7510 Y0.n889 Y0.n888 0.0360676
R7511 Y0.n888 Y0.n887 0.0360676
R7512 Y0.n887 Y0.n274 0.0360676
R7513 Y0.n883 Y0.n274 0.0360676
R7514 Y0.n883 Y0.n882 0.0360676
R7515 Y0.n882 Y0.n881 0.0360676
R7516 Y0.n881 Y0.n279 0.0360676
R7517 Y0.n877 Y0.n279 0.0360676
R7518 Y0.n877 Y0.n876 0.0360676
R7519 Y0.n876 Y0.n875 0.0360676
R7520 Y0.n875 Y0.n8 0.0360676
R7521 Y0.n1364 Y0.n8 0.0360676
R7522 Y0.n1364 Y0.n5 0.0360676
R7523 Y0.n920 Y0.n245 0.0360676
R7524 Y0.n916 Y0.n245 0.0360676
R7525 Y0.n916 Y0.n915 0.0360676
R7526 Y0.n915 Y0.n914 0.0360676
R7527 Y0.n914 Y0.n250 0.0360676
R7528 Y0.n910 Y0.n250 0.0360676
R7529 Y0.n910 Y0.n909 0.0360676
R7530 Y0.n909 Y0.n908 0.0360676
R7531 Y0.n908 Y0.n255 0.0360676
R7532 Y0.n904 Y0.n255 0.0360676
R7533 Y0.n904 Y0.n903 0.0360676
R7534 Y0.n903 Y0.n902 0.0360676
R7535 Y0.n902 Y0.n260 0.0360676
R7536 Y0.n898 Y0.n260 0.0360676
R7537 Y0.n898 Y0.n897 0.0360676
R7538 Y0.n897 Y0.n896 0.0360676
R7539 Y0.n896 Y0.n265 0.0360676
R7540 Y0.n892 Y0.n265 0.0360676
R7541 Y0.n892 Y0.n891 0.0360676
R7542 Y0.n891 Y0.n890 0.0360676
R7543 Y0.n890 Y0.n270 0.0360676
R7544 Y0.n886 Y0.n270 0.0360676
R7545 Y0.n886 Y0.n885 0.0360676
R7546 Y0.n885 Y0.n884 0.0360676
R7547 Y0.n884 Y0.n275 0.0360676
R7548 Y0.n880 Y0.n275 0.0360676
R7549 Y0.n880 Y0.n879 0.0360676
R7550 Y0.n879 Y0.n878 0.0360676
R7551 Y0.n878 Y0.n280 0.0360676
R7552 Y0.n874 Y0.n280 0.0360676
R7553 Y0.n874 Y0.n7 0.0360676
R7554 Y0.n1365 Y0.n7 0.0360676
R7555 Y0.n1366 Y0.n1365 0.0360676
R7556 Y0.n1292 Y0.n45 0.0360676
R7557 Y0 Y0.n1377 0.0245437
R7558 Y0.n100 Y0.n86 0.0234189
R7559 Y0.n962 Y0.n208 0.0234189
R7560 Y0.n964 Y0.n963 0.0234189
R7561 Y0.n1177 Y0.n85 0.0234189
R7562 Y0.n1369 Y0.n1368 0.0233108
R7563 Y0.n244 Y0.n243 0.0233108
R7564 Y0.n922 Y0.n921 0.0233108
R7565 Y0.n1367 Y0.n1 0.0233108
R7566 Y0.n965 Y0.n964 0.0227703
R7567 Y0.n968 Y0.n208 0.0227703
R7568 Y0.n919 Y0.n244 0.0227703
R7569 Y0.n921 Y0.n920 0.0227703
R7570 Y0.n95 Y0.n88 0.0188784
R7571 Y0.n93 Y0.n83 0.0188784
R7572 Y0.n1212 Y0.n1209 0.0188784
R7573 Y0.n1210 Y0.n75 0.0188784
R7574 Y0.n1221 Y0.n77 0.0188784
R7575 Y0.n1235 Y0.n1234 0.0188784
R7576 Y0.n1237 Y0.n64 0.0188784
R7577 Y0.n1249 Y0.n65 0.0188784
R7578 Y0.n1244 Y0.n59 0.0188784
R7579 Y0.n1261 Y0.n1260 0.0188784
R7580 Y0.n1269 Y0.n1268 0.0188784
R7581 Y0.n1274 Y0.n1273 0.0188784
R7582 Y0.n1276 Y0.n47 0.0188784
R7583 Y0.n1289 Y0.n48 0.0188784
R7584 Y0.n1281 Y0.n42 0.0188784
R7585 Y0.n1299 Y0.n1298 0.0188784
R7586 Y0.n1304 Y0.n1303 0.0188784
R7587 Y0.n1307 Y0.n1306 0.0188784
R7588 Y0.n34 Y0.n25 0.0188784
R7589 Y0.n1333 Y0.n1332 0.0188784
R7590 Y0.n1337 Y0.n1336 0.0188784
R7591 Y0.n1341 Y0.n1340 0.0188784
R7592 Y0.n1346 Y0.n1345 0.0188784
R7593 Y0.n469 Y0.n468 0.0188784
R7594 Y0.n477 Y0.n476 0.0188784
R7595 Y0.n486 Y0.n485 0.0188784
R7596 Y0.n495 Y0.n494 0.0188784
R7597 Y0.n502 Y0.n501 0.0188784
R7598 Y0.n528 Y0.n527 0.0188784
R7599 Y0.n536 Y0.n535 0.0188784
R7600 Y0.n543 Y0.n542 0.0188784
R7601 Y0.n558 Y0.n391 0.0188784
R7602 Y0.n561 Y0.n560 0.0188784
R7603 Y0.n575 Y0.n384 0.0188784
R7604 Y0.n585 Y0.n584 0.0188784
R7605 Y0.n594 Y0.n593 0.0188784
R7606 Y0.n603 Y0.n602 0.0188784
R7607 Y0.n612 Y0.n611 0.0188784
R7608 Y0.n619 Y0.n618 0.0188784
R7609 Y0.n630 Y0.n628 0.0188784
R7610 Y0.n644 Y0.n360 0.0188784
R7611 Y0.n660 Y0.n659 0.0188784
R7612 Y0.n675 Y0.n348 0.0188784
R7613 Y0.n678 Y0.n677 0.0188784
R7614 Y0.n686 Y0.n685 0.0188784
R7615 Y0.n701 Y0.n339 0.0188784
R7616 Y0.n445 Y0.n207 0.0188784
R7617 Y0.n971 Y0.n970 0.0188784
R7618 Y0.n980 Y0.n979 0.0188784
R7619 Y0.n982 Y0.n198 0.0188784
R7620 Y0.n1066 Y0.n154 0.0188784
R7621 Y0.n1082 Y0.n1081 0.0188784
R7622 Y0.n1091 Y0.n1090 0.0188784
R7623 Y0.n1093 Y0.n145 0.0188784
R7624 Y0.n727 Y0.n726 0.0188784
R7625 Y0.n736 Y0.n735 0.0188784
R7626 Y0.n740 Y0.n739 0.0188784
R7627 Y0.n744 Y0.n319 0.0188784
R7628 Y0.n805 Y0.n804 0.0188784
R7629 Y0.n809 Y0.n808 0.0188784
R7630 Y0.n816 Y0.n301 0.0188784
R7631 Y0.n819 Y0.n818 0.0188784
R7632 Y0.n1193 Y0.n87 0.0187703
R7633 Y0.n1201 Y0.n88 0.0187703
R7634 Y0.n1229 Y0.n71 0.0187703
R7635 Y0.n1234 Y0.n69 0.0187703
R7636 Y0.n1270 Y0.n1269 0.0187703
R7637 Y0.n1306 Y0.n30 0.0187703
R7638 Y0.n1321 Y0.n31 0.0187703
R7639 Y0.n1347 Y0.n1346 0.0187703
R7640 Y0.n1351 Y0.n1350 0.0187703
R7641 Y0.n453 Y0.n452 0.0187703
R7642 Y0.n468 Y0.n423 0.0187703
R7643 Y0.n513 Y0.n511 0.0187703
R7644 Y0.n527 Y0.n403 0.0187703
R7645 Y0.n576 Y0.n575 0.0187703
R7646 Y0.n645 Y0.n644 0.0187703
R7647 Y0.n653 Y0.n652 0.0187703
R7648 Y0.n702 Y0.n701 0.0187703
R7649 Y0.n711 Y0.n710 0.0187703
R7650 Y0.n996 Y0.n194 0.0187703
R7651 Y0.n1005 Y0.n188 0.0187703
R7652 Y0.n1007 Y0.n185 0.0187703
R7653 Y0.n1013 Y0.n186 0.0187703
R7654 Y0.n1030 Y0.n1029 0.0187703
R7655 Y0.n181 Y0.n179 0.0187703
R7656 Y0.n1040 Y0.n1039 0.0187703
R7657 Y0.n1044 Y0.n1043 0.0187703
R7658 Y0.n1048 Y0.n1047 0.0187703
R7659 Y0.n1053 Y0.n1052 0.0187703
R7660 Y0.n1055 Y0.n158 0.0187703
R7661 Y0.n1071 Y0.n159 0.0187703
R7662 Y0.n1107 Y0.n141 0.0187703
R7663 Y0.n1116 Y0.n135 0.0187703
R7664 Y0.n1118 Y0.n132 0.0187703
R7665 Y0.n1124 Y0.n133 0.0187703
R7666 Y0.n1143 Y0.n1142 0.0187703
R7667 Y0.n1134 Y0.n128 0.0187703
R7668 Y0.n1137 Y0.n1135 0.0187703
R7669 Y0.n1153 Y0.n1152 0.0187703
R7670 Y0.n1155 Y0.n110 0.0187703
R7671 Y0.n1171 Y0.n111 0.0187703
R7672 Y0.n1163 Y0.n106 0.0187703
R7673 Y0.n1183 Y0.n1182 0.0187703
R7674 Y0.n750 Y0.n749 0.0187703
R7675 Y0.n754 Y0.n753 0.0187703
R7676 Y0.n759 Y0.n315 0.0187703
R7677 Y0.n762 Y0.n761 0.0187703
R7678 Y0.n765 Y0.n764 0.0187703
R7679 Y0.n775 Y0.n774 0.0187703
R7680 Y0.n779 Y0.n778 0.0187703
R7681 Y0.n783 Y0.n782 0.0187703
R7682 Y0.n787 Y0.n786 0.0187703
R7683 Y0.n791 Y0.n790 0.0187703
R7684 Y0.n798 Y0.n305 0.0187703
R7685 Y0.n801 Y0.n800 0.0187703
R7686 Y0.n826 Y0.n825 0.0187703
R7687 Y0.n833 Y0.n297 0.0187703
R7688 Y0.n836 Y0.n835 0.0187703
R7689 Y0.n841 Y0.n840 0.0187703
R7690 Y0.n844 Y0.n843 0.0187703
R7691 Y0.n853 Y0.n852 0.0187703
R7692 Y0.n857 Y0.n856 0.0187703
R7693 Y0.n861 Y0.n860 0.0187703
R7694 Y0.n863 Y0.n283 0.0187703
R7695 Y0.n872 Y0.n284 0.0187703
R7696 Y0.n288 Y0.n9 0.0187703
R7697 Y0.n1362 Y0.n11 0.0187703
R7698 Y0.n94 Y0.n93 0.0185541
R7699 Y0.n1341 Y0.n19 0.0185541
R7700 Y0.n476 Y0.n212 0.0185541
R7701 Y0.n685 Y0.n241 0.0185541
R7702 Y0.n988 Y0.n199 0.0184459
R7703 Y0.n1099 Y0.n146 0.0184459
R7704 Y0.n746 Y0.n251 0.0184459
R7705 Y0.n822 Y0.n272 0.0184459
R7706 Y0.n1273 Y0.n53 0.0182297
R7707 Y0.n584 Y0.n226 0.0182297
R7708 Y0.n989 Y0.n988 0.0181216
R7709 Y0.n1100 Y0.n1099 0.0181216
R7710 Y0.n746 Y0.n745 0.0181216
R7711 Y0.n822 Y0.n271 0.0181216
R7712 Y0.n1229 Y0.n1228 0.0175811
R7713 Y0.n1322 Y0.n1321 0.0175811
R7714 Y0.n513 Y0.n512 0.0175811
R7715 Y0.n652 Y0.n235 0.0175811
R7716 Y0.n996 Y0.n995 0.0173649
R7717 Y0.n1107 Y0.n1106 0.0173649
R7718 Y0.n750 Y0.n252 0.0173649
R7719 Y0.n826 Y0.n273 0.0173649
R7720 Y0.n982 Y0.n981 0.0170405
R7721 Y0.n1093 Y0.n1092 0.0170405
R7722 Y0.n319 Y0.n248 0.0170405
R7723 Y0.n818 Y0.n817 0.0170405
R7724 Y0.n1237 Y0.n1236 0.0167162
R7725 Y0.n1305 Y0.n1304 0.0167162
R7726 Y0.n535 Y0.n220 0.0167162
R7727 Y0.n630 Y0.n629 0.0167162
R7728 Y0.n1006 Y0.n1005 0.0162838
R7729 Y0.n1117 Y0.n1116 0.0162838
R7730 Y0.n754 Y0.n253 0.0162838
R7731 Y0.n834 Y0.n833 0.0162838
R7732 Y0.n1260 Y0.n55 0.0159595
R7733 Y0.n1290 Y0.n1289 0.0159595
R7734 Y0.n560 Y0.n225 0.0159595
R7735 Y0.n602 Y0.n373 0.0159595
R7736 Y0.n979 Y0.n201 0.0159595
R7737 Y0.n1090 Y0.n148 0.0159595
R7738 Y0.n739 Y0.n247 0.0159595
R7739 Y0.n301 Y0.n268 0.0159595
R7740 Y0.n1202 Y0.n87 0.0157432
R7741 Y0.n1350 Y0.n3 0.0157432
R7742 Y0.n452 Y0.n211 0.0157432
R7743 Y0.n710 Y0.n242 0.0157432
R7744 Y0.n1209 Y0.n1208 0.0152027
R7745 Y0.n1337 Y0.n21 0.0152027
R7746 Y0.n485 Y0.n416 0.0152027
R7747 Y0.n677 Y0.n240 0.0152027
R7748 Y0.n1014 Y0.n185 0.0152027
R7749 Y0.n1125 Y0.n132 0.0152027
R7750 Y0.n760 Y0.n759 0.0152027
R7751 Y0.n836 Y0.n276 0.0152027
R7752 Y0.n1276 Y0.n1275 0.0148784
R7753 Y0.n593 Y0.n227 0.0148784
R7754 Y0.n970 Y0.n969 0.0148784
R7755 Y0.n1081 Y0.n1080 0.0148784
R7756 Y0.n735 Y0.n246 0.0148784
R7757 Y0.n808 Y0.n267 0.0148784
R7758 Y0.n77 Y0.n76 0.0141216
R7759 Y0.n34 Y0.n33 0.0141216
R7760 Y0.n501 Y0.n217 0.0141216
R7761 Y0.n659 Y0.n236 0.0141216
R7762 Y0.n186 Y0.n178 0.0141216
R7763 Y0.n133 Y0.n126 0.0141216
R7764 Y0.n762 Y0.n256 0.0141216
R7765 Y0.n841 Y0.n277 0.0141216
R7766 Y0.n1178 Y0.n1177 0.0137973
R7767 Y0.n1179 Y0.n100 0.0137973
R7768 Y0.n1066 Y0.n1065 0.0137973
R7769 Y0.n1190 Y0.n99 0.0137973
R7770 Y0.n804 Y0.n266 0.0137973
R7771 Y0.n10 Y0.n6 0.0137973
R7772 Y0.n1368 Y0.n5 0.0137973
R7773 Y0.n1367 Y0.n1366 0.0137973
R7774 Y0.n867 Y0.n15 0.0134381
R7775 Y0.n1250 Y0.n1249 0.0133649
R7776 Y0.n1299 Y0.n40 0.0133649
R7777 Y0.n542 Y0.n221 0.0133649
R7778 Y0.n618 Y0.n232 0.0133649
R7779 Y0.n1029 Y0.n1028 0.0130405
R7780 Y0.n1142 Y0.n1141 0.0130405
R7781 Y0.n764 Y0.n257 0.0130405
R7782 Y0.n843 Y0.n278 0.0130405
R7783 Y0.n1072 Y0.n1071 0.0128243
R7784 Y0.n1183 Y0.n1181 0.0128243
R7785 Y0.n800 Y0.n799 0.0128243
R7786 Y0.n1363 Y0.n1362 0.0128243
R7787 Y0.n1259 Y0.n59 0.0126081
R7788 Y0.n1281 Y0.n1280 0.0126081
R7789 Y0.n559 Y0.n558 0.0126081
R7790 Y0.n611 Y0.n230 0.0126081
R7791 Y0.n1192 Y0.n1191 0.0123919
R7792 Y0.n13 Y0.n4 0.0123919
R7793 Y0.n446 Y0.n210 0.0123919
R7794 Y0.n724 Y0.n332 0.0123919
R7795 Y0.n179 Y0.n171 0.0119595
R7796 Y0.n1138 Y0.n1134 0.0119595
R7797 Y0.n775 Y0.n258 0.0119595
R7798 Y0.n853 Y0.n293 0.0119595
R7799 Y0.n1211 Y0.n1210 0.0118514
R7800 Y0.n1333 Y0.n23 0.0118514
R7801 Y0.n494 Y0.n215 0.0118514
R7802 Y0.n676 Y0.n675 0.0118514
R7803 Y0.n1055 Y0.n1054 0.0117432
R7804 Y0.n1163 Y0.n1162 0.0117432
R7805 Y0.n305 Y0.n263 0.0117432
R7806 Y0.n288 Y0.n287 0.0117432
R7807 Y0.n1188 Y0.n97 0.0116588
R7808 Y0.n1191 Y0.n1190 0.011527
R7809 Y0.n446 Y0.n445 0.011527
R7810 Y0.n13 Y0.n6 0.0114189
R7811 Y0.n727 Y0.n724 0.0114189
R7812 Y0.n325 Y0.n324 0.0109762
R7813 Y0.n323 Y0.n322 0.0109762
R7814 Y0.n768 Y0.n313 0.0109762
R7815 Y0.n771 Y0.n770 0.0109762
R7816 Y0.n769 Y0.n307 0.0109762
R7817 Y0.n795 Y0.n794 0.0109762
R7818 Y0.n812 Y0.n303 0.0109762
R7819 Y0.n813 Y0.n299 0.0109762
R7820 Y0.n830 Y0.n829 0.0109762
R7821 Y0.n847 Y0.n295 0.0109762
R7822 Y0.n849 Y0.n848 0.0109762
R7823 Y0.n866 Y0.n290 0.0109762
R7824 Y0.n868 Y0.n867 0.0109762
R7825 Y0.n1197 Y0.n1196 0.0109762
R7826 Y0.n1197 Y0.n79 0.0109762
R7827 Y0.n1215 Y0.n79 0.0109762
R7828 Y0.n1216 Y0.n1215 0.0109762
R7829 Y0.n1217 Y0.n1216 0.0109762
R7830 Y0.n1217 Y0.n67 0.0109762
R7831 Y0.n1240 Y0.n67 0.0109762
R7832 Y0.n1241 Y0.n1240 0.0109762
R7833 Y0.n1241 Y0.n57 0.0109762
R7834 Y0.n1264 Y0.n57 0.0109762
R7835 Y0.n1265 Y0.n1264 0.0109762
R7836 Y0.n1279 Y0.n51 0.0109762
R7837 Y0.n1286 Y0.n1279 0.0109762
R7838 Y0.n1286 Y0.n1285 0.0109762
R7839 Y0.n1285 Y0.n36 0.0109762
R7840 Y0.n1310 Y0.n36 0.0109762
R7841 Y0.n1311 Y0.n1310 0.0109762
R7842 Y0.n1317 Y0.n1311 0.0109762
R7843 Y0.n1317 Y0.n1316 0.0109762
R7844 Y0.n1316 Y0.n1313 0.0109762
R7845 Y0.n1313 Y0.n1312 0.0109762
R7846 Y0.n1312 Y0.n17 0.0109762
R7847 Y0.n1354 Y0.n17 0.0109762
R7848 Y0.n976 Y0.n192 0.0109762
R7849 Y0.n1002 Y0.n1001 0.0109762
R7850 Y0.n1033 Y0.n175 0.0109762
R7851 Y0.n1036 Y0.n1034 0.0109762
R7852 Y0.n1035 Y0.n163 0.0109762
R7853 Y0.n1061 Y0.n1060 0.0109762
R7854 Y0.n1086 Y0.n152 0.0109762
R7855 Y0.n1087 Y0.n139 0.0109762
R7856 Y0.n1113 Y0.n1112 0.0109762
R7857 Y0.n1146 Y0.n123 0.0109762
R7858 Y0.n1148 Y0.n1147 0.0109762
R7859 Y0.n324 Y0.n323 0.01095
R7860 Y0.n322 Y0.n313 0.01095
R7861 Y0.n771 Y0.n768 0.01095
R7862 Y0.n770 Y0.n769 0.01095
R7863 Y0.n794 Y0.n307 0.01095
R7864 Y0.n795 Y0.n303 0.01095
R7865 Y0.n813 Y0.n812 0.01095
R7866 Y0.n829 Y0.n299 0.01095
R7867 Y0.n830 Y0.n295 0.01095
R7868 Y0.n849 Y0.n847 0.01095
R7869 Y0.n848 Y0.n290 0.01095
R7870 Y0.n868 Y0.n866 0.01095
R7871 Y0.n1265 Y0.n51 0.01095
R7872 Y0.n1355 Y0.n1354 0.01095
R7873 Y0.n976 Y0.n975 0.01095
R7874 Y0.n1001 Y0.n192 0.01095
R7875 Y0.n1002 Y0.n175 0.01095
R7876 Y0.n1034 Y0.n1033 0.01095
R7877 Y0.n1036 Y0.n1035 0.01095
R7878 Y0.n1060 Y0.n163 0.01095
R7879 Y0.n1061 Y0.n152 0.01095
R7880 Y0.n1087 Y0.n1086 0.01095
R7881 Y0.n1112 Y0.n139 0.01095
R7882 Y0.n1113 Y0.n123 0.01095
R7883 Y0.n1147 Y0.n1146 0.01095
R7884 Y0.n1149 Y0.n1148 0.01095
R7885 Y0.n1040 Y0.n169 0.0108784
R7886 Y0.n1135 Y0.n117 0.0108784
R7887 Y0.n779 Y0.n310 0.0108784
R7888 Y0.n857 Y0.n281 0.0108784
R7889 Y0.n1222 Y0.n75 0.0107703
R7890 Y0.n1332 Y0.n1331 0.0107703
R7891 Y0.n495 Y0.n216 0.0107703
R7892 Y0.n348 Y0.n237 0.0107703
R7893 Y0.n1052 Y0.n165 0.0106622
R7894 Y0.n1172 Y0.n1171 0.0106622
R7895 Y0.n790 Y0.n262 0.0106622
R7896 Y0.n873 Y0.n872 0.0106622
R7897 Y0.n1196 Y0.n97 0.0106095
R7898 Y0.n1244 Y0.n1243 0.0100135
R7899 Y0.n1297 Y0.n42 0.0100135
R7900 Y0.n391 Y0.n222 0.0100135
R7901 Y0.n612 Y0.n231 0.0100135
R7902 Y0.n1044 Y0.n167 0.0097973
R7903 Y0.n1154 Y0.n1153 0.0097973
R7904 Y0.n783 Y0.n261 0.0097973
R7905 Y0.n861 Y0.n282 0.0097973
R7906 Y0.n1188 Y0.n1187 0.00967266
R7907 Y0.n1047 Y0.n167 0.00958108
R7908 Y0.n1155 Y0.n1154 0.00958108
R7909 Y0.n786 Y0.n261 0.00958108
R7910 Y0.n863 Y0.n282 0.00958108
R7911 Y0.n1243 Y0.n65 0.00925676
R7912 Y0.n1298 Y0.n1297 0.00925676
R7913 Y0.n543 Y0.n222 0.00925676
R7914 Y0.n619 Y0.n231 0.00925676
R7915 Y0.n1060 Y0.n162 0.00880612
R7916 Y0.n1048 Y0.n165 0.00871622
R7917 Y0.n1172 Y0.n110 0.00871622
R7918 Y0.n787 Y0.n262 0.00871622
R7919 Y0.n873 Y0.n283 0.00871622
R7920 Y0.n1222 Y0.n1221 0.0085
R7921 Y0.n1331 Y0.n25 0.0085
R7922 Y0.n502 Y0.n216 0.0085
R7923 Y0.n660 Y0.n237 0.0085
R7924 Y0.n1043 Y0.n169 0.0085
R7925 Y0.n1152 Y0.n117 0.0085
R7926 Y0.n782 Y0.n310 0.0085
R7927 Y0.n860 Y0.n281 0.0085
R7928 Y0.n326 Y0.n325 0.00809524
R7929 Y0.n1186 Y0.n103 0.00778095
R7930 Y0.n1054 Y0.n1053 0.00763514
R7931 Y0.n1162 Y0.n111 0.00763514
R7932 Y0.n791 Y0.n263 0.00763514
R7933 Y0.n287 Y0.n284 0.00763514
R7934 Y0.n1212 Y0.n1211 0.00741892
R7935 Y0.n1336 Y0.n23 0.00741892
R7936 Y0.n486 Y0.n215 0.00741892
R7937 Y0.n678 Y0.n676 0.00741892
R7938 Y0.n1039 Y0.n171 0.00741892
R7939 Y0.n1138 Y0.n1137 0.00741892
R7940 Y0.n778 Y0.n258 0.00741892
R7941 Y0.n856 Y0.n293 0.00741892
R7942 Y0.n1149 Y0.n115 0.00725714
R7943 Y0.n1187 Y0.n1186 0.00707381
R7944 Y0.n1193 Y0.n1192 0.00698649
R7945 Y0.n1351 Y0.n4 0.00698649
R7946 Y0.n453 Y0.n210 0.00698649
R7947 Y0.n711 Y0.n332 0.00698649
R7948 Y0.n975 Y0.n205 0.00696162
R7949 Y0.n1357 Y0.n1355 0.00691667
R7950 Y0.n1261 Y0.n1259 0.00666216
R7951 Y0.n1280 Y0.n48 0.00666216
R7952 Y0.n561 Y0.n559 0.00666216
R7953 Y0.n603 Y0.n230 0.00666216
R7954 Y0.n1072 Y0.n158 0.00655405
R7955 Y0.n1181 Y0.n106 0.00655405
R7956 Y0.n799 Y0.n798 0.00655405
R7957 Y0.n1363 Y0.n9 0.00655405
R7958 Y0.n1028 Y0.n181 0.00633784
R7959 Y0.n1141 Y0.n128 0.00633784
R7960 Y0.n774 Y0.n257 0.00633784
R7961 Y0.n852 Y0.n278 0.00633784
R7962 Y0.n1250 Y0.n64 0.00590541
R7963 Y0.n1303 Y0.n40 0.00590541
R7964 Y0.n536 Y0.n221 0.00590541
R7965 Y0.n628 Y0.n232 0.00590541
R7966 Y0.n1086 Y0.n151 0.00588776
R7967 Y0.n975 Y0.n204 0.00588776
R7968 Y0.n1065 Y0.n159 0.00547297
R7969 Y0.n1182 Y0.n99 0.00547297
R7970 Y0.n801 Y0.n266 0.00547297
R7971 Y0.n11 Y0.n10 0.00547297
R7972 Y0.n1030 Y0.n178 0.00525676
R7973 Y0.n1143 Y0.n126 0.00525676
R7974 Y0.n765 Y0.n256 0.00525676
R7975 Y0.n844 Y0.n277 0.00525676
R7976 Y0.n76 Y0.n71 0.00514865
R7977 Y0.n33 Y0.n31 0.00514865
R7978 Y0.n511 Y0.n217 0.00514865
R7979 Y0.n653 Y0.n236 0.00514865
R7980 Y0.n1356 Y0.n15 0.00440238
R7981 Y0.n1275 Y0.n1274 0.00439189
R7982 Y0.n585 Y0.n227 0.00439189
R7983 Y0.n969 Y0.n207 0.00439189
R7984 Y0.n1080 Y0.n154 0.00439189
R7985 Y0.n726 Y0.n246 0.00439189
R7986 Y0.n805 Y0.n267 0.00439189
R7987 Y0.n1194 Y0.n98 0.00425921
R7988 Y0.n1200 Y0.n89 0.00425921
R7989 Y0.n82 Y0.n81 0.00425921
R7990 Y0.n1220 Y0.n1219 0.00425921
R7991 Y0.n1233 Y0.n68 0.00425921
R7992 Y0.n1238 Y0.n66 0.00425921
R7993 Y0.n1248 Y0.n1247 0.00425921
R7994 Y0.n1245 Y0.n58 0.00425921
R7995 Y0.n1272 Y0.n52 0.00425921
R7996 Y0.n1283 Y0.n1282 0.00425921
R7997 Y0.n1300 Y0.n41 0.00425921
R7998 Y0.n1302 Y0.n37 0.00425921
R7999 Y0.n1308 Y0.n39 0.00425921
R8000 Y0.n1314 Y0.n35 0.00425921
R8001 Y0.n1334 Y0.n24 0.00425921
R8002 Y0.n1349 Y0.n1348 0.00425921
R8003 Y0.n1352 Y0.n14 0.00425921
R8004 Y0.n1042 Y0.n1041 0.00425921
R8005 Y0.n1046 Y0.n1045 0.00425921
R8006 Y0.n1151 Y0.n118 0.00425921
R8007 Y0.n1156 Y0.n116 0.00425921
R8008 Y0.n743 Y0.n742 0.00425921
R8009 Y0.n748 Y0.n747 0.00425921
R8010 Y0.n752 Y0.n751 0.00425921
R8011 Y0.n756 Y0.n755 0.00425921
R8012 Y0.n777 Y0.n776 0.00425921
R8013 Y0.n781 Y0.n780 0.00425921
R8014 Y0.n785 Y0.n784 0.00425921
R8015 Y0.n789 Y0.n788 0.00425921
R8016 Y0.n806 Y0.n803 0.00425921
R8017 Y0.n820 Y0.n300 0.00425921
R8018 Y0.n824 Y0.n823 0.00425921
R8019 Y0.n827 Y0.n298 0.00425921
R8020 Y0.n832 Y0.n296 0.00425921
R8021 Y0.n855 Y0.n854 0.00425921
R8022 Y0.n859 Y0.n858 0.00425921
R8023 Y0.n864 Y0.n862 0.00425921
R8024 Y0.n871 Y0.n285 0.00425921
R8025 Y0.n1161 Y0.n1160 0.00424524
R8026 Y0.n1200 Y0.n1199 0.0042371
R8027 Y0.n96 Y0.n92 0.0042371
R8028 Y0.n90 Y0.n80 0.0042371
R8029 Y0.n1213 Y0.n82 0.0042371
R8030 Y0.n1230 Y0.n70 0.0042371
R8031 Y0.n1233 Y0.n1232 0.0042371
R8032 Y0.n1262 Y0.n58 0.0042371
R8033 Y0.n1267 Y0.n56 0.0042371
R8034 Y0.n1271 Y0.n54 0.0042371
R8035 Y0.n1272 Y0.n1271 0.0042371
R8036 Y0.n1277 Y0.n52 0.0042371
R8037 Y0.n1288 Y0.n49 0.0042371
R8038 Y0.n1282 Y0.n50 0.0042371
R8039 Y0.n39 Y0.n38 0.0042371
R8040 Y0.n1320 Y0.n1319 0.0042371
R8041 Y0.n1335 Y0.n1334 0.0042371
R8042 Y0.n1339 Y0.n1338 0.0042371
R8043 Y0.n1344 Y0.n1342 0.0042371
R8044 Y0.n1348 Y0.n18 0.0042371
R8045 Y0.n983 Y0.n200 0.0042371
R8046 Y0.n1012 Y0.n176 0.0042371
R8047 Y0.n1031 Y0.n177 0.0042371
R8048 Y0.n1070 Y0.n1069 0.0042371
R8049 Y0.n1094 Y0.n147 0.0042371
R8050 Y0.n1123 Y0.n124 0.0042371
R8051 Y0.n1144 Y0.n125 0.0042371
R8052 Y0.n1164 Y0.n104 0.0042371
R8053 Y0.n1184 Y0.n105 0.0042371
R8054 Y0.n738 Y0.n737 0.0042371
R8055 Y0.n742 Y0.n741 0.0042371
R8056 Y0.n758 Y0.n756 0.0042371
R8057 Y0.n763 Y0.n314 0.0042371
R8058 Y0.n766 Y0.n312 0.0042371
R8059 Y0.n776 Y0.n773 0.0042371
R8060 Y0.n792 Y0.n789 0.0042371
R8061 Y0.n797 Y0.n306 0.0042371
R8062 Y0.n802 Y0.n304 0.0042371
R8063 Y0.n803 Y0.n802 0.0042371
R8064 Y0.n807 Y0.n806 0.0042371
R8065 Y0.n810 Y0.n302 0.0042371
R8066 Y0.n815 Y0.n300 0.0042371
R8067 Y0.n837 Y0.n296 0.0042371
R8068 Y0.n842 Y0.n839 0.0042371
R8069 Y0.n845 Y0.n294 0.0042371
R8070 Y0.n854 Y0.n851 0.0042371
R8071 Y0.n871 Y0.n870 0.0042371
R8072 Y0.n289 Y0.n286 0.0042371
R8073 Y0.n1361 Y0.n1360 0.0042371
R8074 Y0.n1360 Y0.n1359 0.0042371
R8075 Y0.n730 Y0.n729 0.00423273
R8076 Y0.n441 Y0.n440 0.00422178
R8077 Y0.n717 Y0.n329 0.00422178
R8078 Y0.n1159 Y0.n115 0.00421905
R8079 Y0.n1014 Y0.n1013 0.00417568
R8080 Y0.n1125 Y0.n1124 0.00417568
R8081 Y0.n761 Y0.n760 0.00417568
R8082 Y0.n840 Y0.n276 0.00417568
R8083 Y0.n1198 Y0.n96 0.00410442
R8084 Y0.n1344 Y0.n1343 0.00410442
R8085 Y0.n1208 Y0.n83 0.00406757
R8086 Y0.n1340 Y0.n21 0.00406757
R8087 Y0.n477 Y0.n416 0.00406757
R8088 Y0.n686 Y0.n240 0.00406757
R8089 Y0.n1056 Y0.n160 0.00402269
R8090 Y0.n987 Y0.n190 0.00398793
R8091 Y0.n1098 Y0.n137 0.00398793
R8092 Y0.n747 Y0.n318 0.00397174
R8093 Y0.n785 Y0.n308 0.00397174
R8094 Y0.n823 Y0.n821 0.00397174
R8095 Y0.n865 Y0.n864 0.00397174
R8096 Y0.n1247 Y0.n1246 0.00394963
R8097 Y0.n1284 Y0.n41 0.00394963
R8098 Y0.n978 Y0.n202 0.00394626
R8099 Y0.n1089 Y0.n149 0.00394626
R8100 Y0.n433 Y0.n203 0.00393696
R8101 Y0.n1063 Y0.n150 0.00393696
R8102 Y0.n997 Y0.n189 0.00390294
R8103 Y0.n1108 Y0.n136 0.00390294
R8104 Y0.n1051 Y0.n161 0.00389381
R8105 Y0.n1008 Y0.n187 0.00385851
R8106 Y0.n1037 Y0.n172 0.00385851
R8107 Y0.n1119 Y0.n134 0.00385851
R8108 Y0.n1133 Y0.n119 0.00385851
R8109 Y0.n1009 Y0.n1008 0.00380768
R8110 Y0.n1120 Y0.n1119 0.00380768
R8111 Y0.n174 Y0.n172 0.00380053
R8112 Y0.n1133 Y0.n122 0.00380053
R8113 Y0.n1220 Y0.n78 0.00379484
R8114 Y0.n1315 Y0.n1314 0.00379484
R8115 Y0.n728 Y0.n328 0.00379484
R8116 Y0.n1189 Y0.n102 0.00377273
R8117 Y0.n984 Y0.n983 0.0037725
R8118 Y0.n1051 Y0.n1050 0.0037725
R8119 Y0.n1095 Y0.n1094 0.0037725
R8120 Y0.n1168 Y0.n1167 0.00374762
R8121 Y0.n1064 Y0.n1063 0.00372958
R8122 Y0.n757 Y0.n314 0.0037285
R8123 Y0.n839 Y0.n838 0.0037285
R8124 Y0.n1069 Y0.n1068 0.00372177
R8125 Y0.n772 Y0.n312 0.00370639
R8126 Y0.n850 Y0.n294 0.00370639
R8127 Y0.n1166 Y0.n103 0.00369524
R8128 Y0.n1231 Y0.n1230 0.00366216
R8129 Y0.n1320 Y0.n32 0.00366216
R8130 Y0.n114 Y0.n112 0.00366216
R8131 Y0.n1158 Y0.n1157 0.00364005
R8132 Y0.n1202 Y0.n1201 0.00363514
R8133 Y0.n1347 Y0.n3 0.00363514
R8134 Y0.n423 Y0.n211 0.00363514
R8135 Y0.n702 Y0.n242 0.00363514
R8136 Y0.n733 Y0.n731 0.00359048
R8137 Y0.n1046 Y0.n166 0.00358532
R8138 Y0.n440 Y0.n436 0.00357902
R8139 Y0.n717 Y0.n716 0.00357902
R8140 Y0.n987 Y0.n986 0.00357098
R8141 Y0.n1098 Y0.n1097 0.00357098
R8142 Y0.n1239 Y0.n1238 0.00348526
R8143 Y0.n1309 Y0.n37 0.00348526
R8144 Y0.n1012 Y0.n1011 0.003457
R8145 Y0.n1123 Y0.n1122 0.003457
R8146 Y0.n177 Y0.n173 0.00344926
R8147 Y0.n125 Y0.n121 0.00344926
R8148 Y0.n752 Y0.n316 0.00344103
R8149 Y0.n780 Y0.n311 0.00344103
R8150 Y0.n831 Y0.n298 0.00344103
R8151 Y0.n858 Y0.n292 0.00344103
R8152 Y0.n1038 Y0.n170 0.00343273
R8153 Y0.n1136 Y0.n120 0.00343273
R8154 Y0.n1004 Y0.n1003 0.00341839
R8155 Y0.n1115 Y0.n1114 0.00341839
R8156 Y0.n1112 Y0.n138 0.00341837
R8157 Y0.n1001 Y0.n191 0.00341837
R8158 Y0.n732 Y0.n326 0.00335476
R8159 Y0.n1214 Y0.n80 0.00335258
R8160 Y0.n1338 Y0.n22 0.00335258
R8161 Y0.n1003 Y0.n189 0.0033136
R8162 Y0.n1114 Y0.n136 0.0033136
R8163 Y0.n1268 Y0.n55 0.00331081
R8164 Y0.n1290 Y0.n47 0.00331081
R8165 Y0.n384 Y0.n225 0.00331081
R8166 Y0.n594 Y0.n373 0.00331081
R8167 Y0.n971 Y0.n201 0.00331081
R8168 Y0.n1082 Y0.n148 0.00331081
R8169 Y0.n736 Y0.n247 0.00331081
R8170 Y0.n809 Y0.n268 0.00331081
R8171 Y0.n180 Y0.n173 0.00330444
R8172 Y0.n127 Y0.n121 0.00330444
R8173 Y0.n1041 Y0.n170 0.0032992
R8174 Y0.n120 Y0.n118 0.0032992
R8175 Y0.n1011 Y0.n1010 0.00329663
R8176 Y0.n1122 Y0.n1121 0.00329663
R8177 Y0.n1169 Y0.n113 0.00324201
R8178 Y0.n1263 Y0.n56 0.00319779
R8179 Y0.n1288 Y0.n1287 0.00319779
R8180 Y0.n1165 Y0.n1164 0.00319779
R8181 Y0.n793 Y0.n306 0.00319779
R8182 Y0.n869 Y0.n289 0.00319779
R8183 Y0.n978 Y0.n977 0.00317568
R8184 Y0.n1089 Y0.n1088 0.00317568
R8185 Y0.n738 Y0.n320 0.00317568
R8186 Y0.n814 Y0.n302 0.00317568
R8187 Y0.n986 Y0.n985 0.00316007
R8188 Y0.n1097 Y0.n1096 0.00316007
R8189 Y0.n1049 Y0.n166 0.00314581
R8190 Y0.n734 Y0.n327 0.00310934
R8191 Y0.n1007 Y0.n1006 0.00309459
R8192 Y0.n1118 Y0.n1117 0.00309459
R8193 Y0.n315 Y0.n253 0.00309459
R8194 Y0.n835 Y0.n834 0.00309459
R8195 Y0.n1195 Y0.n1194 0.003043
R8196 Y0.n1353 Y0.n1352 0.003043
R8197 Y0.n1067 Y0.n1064 0.00302306
R8198 Y0.n1068 Y0.n1067 0.00300884
R8199 Y0.n482 Y0.n480 0.0029881
R8200 Y0.n517 Y0.n516 0.0029881
R8201 Y0.n532 Y0.n398 0.0029881
R8202 Y0.n634 Y0.n633 0.0029881
R8203 Y0.n1050 Y0.n1049 0.00298054
R8204 Y0.n985 Y0.n984 0.00298054
R8205 Y0.n1096 Y0.n1095 0.00298054
R8206 Y0.n649 Y0.n355 0.0029619
R8207 Y0.n683 Y0.n682 0.0029619
R8208 Y0.n180 Y0.n174 0.00293083
R8209 Y0.n127 Y0.n122 0.00293083
R8210 Y0.n1010 Y0.n1009 0.0029237
R8211 Y0.n1121 Y0.n1120 0.0029237
R8212 Y0.n1267 Y0.n1266 0.00291032
R8213 Y0.n1278 Y0.n49 0.00291032
R8214 Y0.n1062 Y0.n160 0.00291032
R8215 Y0.n1185 Y0.n104 0.00291032
R8216 Y0.n737 Y0.n321 0.00291032
R8217 Y0.n797 Y0.n796 0.00291032
R8218 Y0.n811 Y0.n810 0.00291032
R8219 Y0.n286 Y0.n12 0.00291032
R8220 Y0.n1004 Y0.n187 0.00289527
R8221 Y0.n1115 Y0.n134 0.00289527
R8222 Y0.n1038 Y0.n1037 0.00289527
R8223 Y0.n1136 Y0.n119 0.00289527
R8224 Y0.n438 Y0.n436 0.00287188
R8225 Y0.n719 Y0.n716 0.00284569
R8226 Y0.n164 Y0.n161 0.00283826
R8227 Y0.n1357 Y0.n1356 0.00283095
R8228 Y0.n206 Y0.n203 0.00279542
R8229 Y0.n153 Y0.n150 0.00279542
R8230 Y0.n193 Y0.n190 0.00276679
R8231 Y0.n140 Y0.n137 0.00276679
R8232 Y0.n91 Y0.n90 0.00275553
R8233 Y0.n1339 Y0.n20 0.00275553
R8234 Y0.n101 Y0.n98 0.00273342
R8235 Y0.n1359 Y0.n14 0.00273342
R8236 Y0.n438 Y0.n437 0.00272619
R8237 Y0.n437 Y0.n430 0.00272619
R8238 Y0.n456 Y0.n428 0.00272619
R8239 Y0.n458 Y0.n457 0.00272619
R8240 Y0.n466 Y0.n465 0.00272619
R8241 Y0.n474 Y0.n418 0.00272619
R8242 Y0.n479 Y0.n418 0.00272619
R8243 Y0.n481 Y0.n414 0.00272619
R8244 Y0.n489 Y0.n414 0.00272619
R8245 Y0.n497 Y0.n411 0.00272619
R8246 Y0.n498 Y0.n497 0.00272619
R8247 Y0.n507 Y0.n506 0.00272619
R8248 Y0.n508 Y0.n507 0.00272619
R8249 Y0.n518 Y0.n405 0.00272619
R8250 Y0.n522 Y0.n405 0.00272619
R8251 Y0.n530 Y0.n401 0.00272619
R8252 Y0.n531 Y0.n530 0.00272619
R8253 Y0.n539 Y0.n538 0.00272619
R8254 Y0.n540 Y0.n395 0.00272619
R8255 Y0.n552 Y0.n393 0.00272619
R8256 Y0.n564 Y0.n389 0.00272619
R8257 Y0.n565 Y0.n564 0.00272619
R8258 Y0.n571 Y0.n570 0.00272619
R8259 Y0.n573 Y0.n571 0.00272619
R8260 Y0.n573 Y0.n572 0.00272619
R8261 Y0.n582 Y0.n581 0.00272619
R8262 Y0.n591 Y0.n590 0.00272619
R8263 Y0.n590 Y0.n375 0.00272619
R8264 Y0.n600 Y0.n599 0.00272619
R8265 Y0.n599 Y0.n371 0.00272619
R8266 Y0.n606 Y0.n371 0.00272619
R8267 Y0.n614 Y0.n368 0.00272619
R8268 Y0.n615 Y0.n614 0.00272619
R8269 Y0.n624 Y0.n623 0.00272619
R8270 Y0.n625 Y0.n624 0.00272619
R8271 Y0.n639 Y0.n362 0.00272619
R8272 Y0.n648 Y0.n647 0.00272619
R8273 Y0.n656 Y0.n655 0.00272619
R8274 Y0.n657 Y0.n352 0.00272619
R8275 Y0.n669 Y0.n350 0.00272619
R8276 Y0.n681 Y0.n346 0.00272619
R8277 Y0.n682 Y0.n681 0.00272619
R8278 Y0.n689 Y0.n344 0.00272619
R8279 Y0.n690 Y0.n689 0.00272619
R8280 Y0.n691 Y0.n690 0.00272619
R8281 Y0.n699 Y0.n697 0.00272619
R8282 Y0.n699 Y0.n698 0.00272619
R8283 Y0.n708 Y0.n706 0.00272619
R8284 Y0.n708 Y0.n707 0.00272619
R8285 Y0.n722 Y0.n721 0.00272619
R8286 Y0.n720 Y0.n719 0.00272619
R8287 Y0.n448 Y0.n430 0.0027
R8288 Y0.n457 Y0.n456 0.0027
R8289 Y0.n466 Y0.n464 0.0027
R8290 Y0.n474 Y0.n473 0.0027
R8291 Y0.n482 Y0.n481 0.0027
R8292 Y0.n508 Y0.n407 0.0027
R8293 Y0.n540 Y0.n539 0.0027
R8294 Y0.n548 Y0.n393 0.0027
R8295 Y0.n554 Y0.n389 0.0027
R8296 Y0.n582 Y0.n580 0.0027
R8297 Y0.n591 Y0.n589 0.0027
R8298 Y0.n625 Y0.n364 0.0027
R8299 Y0.n635 Y0.n362 0.0027
R8300 Y0.n647 Y0.n358 0.0027
R8301 Y0.n657 Y0.n656 0.0027
R8302 Y0.n665 Y0.n350 0.0027
R8303 Y0.n671 Y0.n346 0.0027
R8304 Y0.n707 Y0.n334 0.0027
R8305 Y0.n721 Y0.n720 0.0027
R8306 Y0.n516 Y0.n407 0.00264762
R8307 Y0.n655 Y0.n355 0.00264762
R8308 Y0.n751 Y0.n317 0.00264496
R8309 Y0.n828 Y0.n827 0.00264496
R8310 Y0.n1042 Y0.n168 0.00262285
R8311 Y0.n1151 Y0.n1150 0.00262285
R8312 Y0.n781 Y0.n309 0.00262285
R8313 Y0.n859 Y0.n291 0.00262285
R8314 Y0.n532 Y0.n531 0.00262143
R8315 Y0.n635 Y0.n634 0.00262143
R8316 Y0.n1242 Y0.n66 0.00260074
R8317 Y0.n1302 Y0.n1301 0.00260074
R8318 Y0.n484 Y0.n417 0.00257862
R8319 Y0.n684 Y0.n345 0.00257862
R8320 Y0.n633 Y0.n364 0.00256905
R8321 Y0.n1236 Y0.n1235 0.00255405
R8322 Y0.n1307 Y0.n1305 0.00255405
R8323 Y0.n528 Y0.n220 0.00255405
R8324 Y0.n629 Y0.n360 0.00255405
R8325 Y0.n538 Y0.n398 0.00254286
R8326 Y0.n649 Y0.n648 0.00254286
R8327 Y0.n534 Y0.n399 0.0025344
R8328 Y0.n518 Y0.n517 0.00251667
R8329 Y0.n632 Y0.n631 0.00251228
R8330 Y0.n443 Y0.n442 0.0024936
R8331 Y0.n480 Y0.n479 0.00246429
R8332 Y0.n683 Y0.n344 0.00246429
R8333 Y0.n1218 Y0.n70 0.00244595
R8334 Y0.n1319 Y0.n1318 0.00244595
R8335 Y0.n499 Y0.n498 0.0024381
R8336 Y0.n665 Y0.n664 0.0024381
R8337 Y0.n515 Y0.n514 0.00242383
R8338 Y0.n651 Y0.n356 0.00242383
R8339 Y0.n731 Y0.n730 0.00238571
R8340 Y0.n1168 Y0.n1161 0.00238571
R8341 Y0.n463 Y0.n426 0.00238571
R8342 Y0.n472 Y0.n421 0.00238571
R8343 Y0.n491 Y0.n490 0.00238571
R8344 Y0.n499 Y0.n409 0.00238571
R8345 Y0.n524 Y0.n523 0.00238571
R8346 Y0.n547 Y0.n546 0.00238571
R8347 Y0.n555 Y0.n553 0.00238571
R8348 Y0.n579 Y0.n382 0.00238571
R8349 Y0.n588 Y0.n378 0.00238571
R8350 Y0.n597 Y0.n375 0.00238571
R8351 Y0.n608 Y0.n607 0.00238571
R8352 Y0.n616 Y0.n366 0.00238571
R8353 Y0.n641 Y0.n640 0.00238571
R8354 Y0.n664 Y0.n663 0.00238571
R8355 Y0.n672 Y0.n670 0.00238571
R8356 Y0.n696 Y0.n342 0.00238571
R8357 Y0.n705 Y0.n337 0.00238571
R8358 Y0.n455 Y0.n454 0.00237961
R8359 Y0.n459 Y0.n427 0.00237961
R8360 Y0.n467 Y0.n425 0.00237961
R8361 Y0.n475 Y0.n419 0.00237961
R8362 Y0.n478 Y0.n419 0.00237961
R8363 Y0.n487 Y0.n415 0.00237961
R8364 Y0.n488 Y0.n487 0.00237961
R8365 Y0.n496 Y0.n412 0.00237961
R8366 Y0.n496 Y0.n410 0.00237961
R8367 Y0.n505 Y0.n408 0.00237961
R8368 Y0.n509 Y0.n408 0.00237961
R8369 Y0.n520 Y0.n519 0.00237961
R8370 Y0.n521 Y0.n520 0.00237961
R8371 Y0.n529 Y0.n402 0.00237961
R8372 Y0.n529 Y0.n400 0.00237961
R8373 Y0.n537 Y0.n397 0.00237961
R8374 Y0.n541 Y0.n396 0.00237961
R8375 Y0.n551 Y0.n550 0.00237961
R8376 Y0.n563 Y0.n562 0.00237961
R8377 Y0.n563 Y0.n388 0.00237961
R8378 Y0.n569 Y0.n385 0.00237961
R8379 Y0.n574 Y0.n385 0.00237961
R8380 Y0.n574 Y0.n386 0.00237961
R8381 Y0.n583 Y0.n381 0.00237961
R8382 Y0.n592 Y0.n376 0.00237961
R8383 Y0.n595 Y0.n376 0.00237961
R8384 Y0.n601 Y0.n372 0.00237961
R8385 Y0.n604 Y0.n372 0.00237961
R8386 Y0.n605 Y0.n604 0.00237961
R8387 Y0.n613 Y0.n369 0.00237961
R8388 Y0.n613 Y0.n367 0.00237961
R8389 Y0.n622 Y0.n365 0.00237961
R8390 Y0.n626 Y0.n365 0.00237961
R8391 Y0.n638 Y0.n637 0.00237961
R8392 Y0.n646 Y0.n357 0.00237961
R8393 Y0.n654 Y0.n354 0.00237961
R8394 Y0.n658 Y0.n353 0.00237961
R8395 Y0.n668 Y0.n667 0.00237961
R8396 Y0.n680 Y0.n679 0.00237961
R8397 Y0.n680 Y0.n345 0.00237961
R8398 Y0.n688 Y0.n687 0.00237961
R8399 Y0.n688 Y0.n343 0.00237961
R8400 Y0.n692 Y0.n343 0.00237961
R8401 Y0.n700 Y0.n340 0.00237961
R8402 Y0.n700 Y0.n341 0.00237961
R8403 Y0.n709 Y0.n336 0.00237961
R8404 Y0.n709 Y0.n335 0.00237961
R8405 Y0.n723 Y0.n330 0.00237961
R8406 Y0.n444 Y0.n435 0.00237961
R8407 Y0.n973 Y0.n972 0.00237961
R8408 Y0.n1032 Y0.n176 0.00237961
R8409 Y0.n1032 Y0.n1031 0.00237961
R8410 Y0.n1058 Y0.n1057 0.00237961
R8411 Y0.n1084 Y0.n1083 0.00237961
R8412 Y0.n1145 Y0.n124 0.00237961
R8413 Y0.n1145 Y0.n1144 0.00237961
R8414 Y0.n767 Y0.n763 0.00237961
R8415 Y0.n767 Y0.n766 0.00237961
R8416 Y0.n846 Y0.n842 0.00237961
R8417 Y0.n846 Y0.n845 0.00237961
R8418 Y0.n548 Y0.n547 0.00235952
R8419 Y0.n570 Y0.n387 0.00235952
R8420 Y0.n447 Y0.n431 0.00235749
R8421 Y0.n455 Y0.n427 0.00235749
R8422 Y0.n467 Y0.n424 0.00235749
R8423 Y0.n475 Y0.n420 0.00235749
R8424 Y0.n483 Y0.n415 0.00235749
R8425 Y0.n510 Y0.n509 0.00235749
R8426 Y0.n541 Y0.n397 0.00235749
R8427 Y0.n550 Y0.n549 0.00235749
R8428 Y0.n562 Y0.n390 0.00235749
R8429 Y0.n583 Y0.n380 0.00235749
R8430 Y0.n592 Y0.n377 0.00235749
R8431 Y0.n627 Y0.n626 0.00235749
R8432 Y0.n637 Y0.n636 0.00235749
R8433 Y0.n646 Y0.n359 0.00235749
R8434 Y0.n658 Y0.n354 0.00235749
R8435 Y0.n667 Y0.n666 0.00235749
R8436 Y0.n679 Y0.n347 0.00235749
R8437 Y0.n712 Y0.n335 0.00235749
R8438 Y0.n999 Y0.n998 0.00235749
R8439 Y0.n1110 Y0.n1109 0.00235749
R8440 Y0.n1372 Y0.n0 0.00233784
R8441 Y0.n616 Y0.n615 0.00233333
R8442 Y0.n515 Y0.n510 0.00231327
R8443 Y0.n654 Y0.n356 0.00231327
R8444 Y0.n449 Y0.n448 0.00230714
R8445 Y0.n714 Y0.n334 0.00230714
R8446 Y0.n722 Y0.n715 0.00230714
R8447 Y0.n1219 Y0.n1218 0.00229115
R8448 Y0.n1318 Y0.n35 0.00229115
R8449 Y0.n533 Y0.n400 0.00229115
R8450 Y0.n636 Y0.n363 0.00229115
R8451 Y0.n450 Y0.n428 0.00228095
R8452 Y0.n465 Y0.n421 0.00228095
R8453 Y0.n697 Y0.n696 0.00225476
R8454 Y0.n632 Y0.n627 0.00224693
R8455 Y0.n981 Y0.n980 0.00222973
R8456 Y0.n1092 Y0.n1091 0.00222973
R8457 Y0.n740 Y0.n248 0.00222973
R8458 Y0.n817 Y0.n816 0.00222973
R8459 Y0.n537 Y0.n399 0.00222482
R8460 Y0.n650 Y0.n357 0.00222482
R8461 Y0.n519 Y0.n406 0.0022027
R8462 Y0.n566 Y0.n565 0.00220238
R8463 Y0.n600 Y0.n598 0.00220238
R8464 Y0.n580 Y0.n579 0.00217619
R8465 Y0.n581 Y0.n378 0.00217619
R8466 Y0.n478 Y0.n417 0.00215848
R8467 Y0.n687 Y0.n684 0.00215848
R8468 Y0.n1248 Y0.n1242 0.00213636
R8469 Y0.n1301 Y0.n1300 0.00213636
R8470 Y0.n500 Y0.n410 0.00213636
R8471 Y0.n666 Y0.n351 0.00213636
R8472 Y0.n1045 Y0.n168 0.00211425
R8473 Y0.n1150 Y0.n116 0.00211425
R8474 Y0.n784 Y0.n309 0.00211425
R8475 Y0.n862 Y0.n291 0.00211425
R8476 Y0.n733 Y0.n732 0.00209762
R8477 Y0.n464 Y0.n463 0.00209762
R8478 Y0.n596 Y0.n595 0.00209214
R8479 Y0.n1000 Y0.n193 0.00209214
R8480 Y0.n1111 Y0.n140 0.00209214
R8481 Y0.n748 Y0.n317 0.00209214
R8482 Y0.n828 Y0.n824 0.00209214
R8483 Y0.n698 Y0.n337 0.00207143
R8484 Y0.n549 Y0.n394 0.00207002
R8485 Y0.n569 Y0.n568 0.00207002
R8486 Y0.n617 Y0.n367 0.00204791
R8487 Y0.n447 Y0.n429 0.0020258
R8488 Y0.n713 Y0.n712 0.0020258
R8489 Y0.n723 Y0.n333 0.0020258
R8490 Y0.n553 Y0.n552 0.00201905
R8491 Y0.n995 Y0.n188 0.00201351
R8492 Y0.n1106 Y0.n135 0.00201351
R8493 Y0.n753 Y0.n252 0.00201351
R8494 Y0.n297 Y0.n273 0.00201351
R8495 Y0.n92 Y0.n91 0.00200369
R8496 Y0.n1342 Y0.n20 0.00200369
R8497 Y0.n454 Y0.n451 0.00200369
R8498 Y0.n425 Y0.n422 0.00200369
R8499 Y0.n443 Y0.n441 0.00200107
R8500 Y0.n442 Y0.n205 0.00200107
R8501 Y0.n729 Y0.n329 0.00200107
R8502 Y0.n608 Y0.n368 0.00199286
R8503 Y0.n695 Y0.n340 0.00198157
R8504 Y0.n567 Y0.n388 0.00193735
R8505 Y0.n601 Y0.n374 0.00193735
R8506 Y0.n578 Y0.n380 0.00191523
R8507 Y0.n381 Y0.n379 0.00191523
R8508 Y0.n444 Y0.n432 0.00191523
R8509 Y0.n435 Y0.n434 0.00191523
R8510 Y0.n728 Y0.n331 0.00191523
R8511 Y0.n1359 Y0.n1358 0.00191523
R8512 Y0.n491 Y0.n411 0.00191429
R8513 Y0.n670 Y0.n669 0.00191429
R8514 Y0.n504 Y0.n503 0.00187101
R8515 Y0.n998 Y0.n997 0.00185493
R8516 Y0.n1109 Y0.n1108 0.00185493
R8517 Y0.n1266 Y0.n54 0.00184889
R8518 Y0.n1278 Y0.n1277 0.00184889
R8519 Y0.n462 Y0.n424 0.00184889
R8520 Y0.n662 Y0.n661 0.00184889
R8521 Y0.n974 Y0.n206 0.00184889
R8522 Y0.n1070 Y0.n1062 0.00184889
R8523 Y0.n1085 Y0.n153 0.00184889
R8524 Y0.n1185 Y0.n1184 0.00184889
R8525 Y0.n734 Y0.n321 0.00184889
R8526 Y0.n796 Y0.n304 0.00184889
R8527 Y0.n811 Y0.n807 0.00184889
R8528 Y0.n1361 Y0.n12 0.00184889
R8529 Y0.n641 Y0.n358 0.00183571
R8530 Y0.n341 Y0.n338 0.00182678
R8531 Y0.n523 Y0.n522 0.00180952
R8532 Y0.n1228 Y0.n69 0.0017973
R8533 Y0.n1322 Y0.n30 0.0017973
R8534 Y0.n512 Y0.n403 0.0017973
R8535 Y0.n645 Y0.n235 0.0017973
R8536 Y0.n972 Y0.n202 0.0017897
R8537 Y0.n1083 Y0.n149 0.0017897
R8538 Y0.n545 Y0.n544 0.00178256
R8539 Y0.n551 Y0.n392 0.00178256
R8540 Y0.n621 Y0.n620 0.00178256
R8541 Y0.n609 Y0.n369 0.00176044
R8542 Y0.n1167 Y0.n1166 0.00175714
R8543 Y0.n524 Y0.n401 0.00173095
R8544 Y0.n640 Y0.n639 0.00173095
R8545 Y0.n471 Y0.n470 0.00171622
R8546 Y0.n1057 Y0.n1056 0.00171347
R8547 Y0.n1195 Y0.n89 0.0016941
R8548 Y0.n1353 Y0.n1349 0.0016941
R8549 Y0.n492 Y0.n412 0.0016941
R8550 Y0.n668 Y0.n349 0.0016941
R8551 Y0.n694 Y0.n693 0.0016941
R8552 Y0.n672 Y0.n671 0.00165238
R8553 Y0.n577 Y0.n383 0.00162776
R8554 Y0.n587 Y0.n586 0.00162776
R8555 Y0.n642 Y0.n359 0.00162776
R8556 Y0.n725 Y0.n327 0.00162776
R8557 Y0.n490 Y0.n489 0.00162619
R8558 Y0.n521 Y0.n404 0.00160565
R8559 Y0.n977 Y0.n200 0.00158354
R8560 Y0.n1088 Y0.n147 0.00158354
R8561 Y0.n741 Y0.n320 0.00158354
R8562 Y0.n815 Y0.n814 0.00158354
R8563 Y0.n1263 Y0.n1262 0.00156143
R8564 Y0.n1287 Y0.n50 0.00156143
R8565 Y0.n461 Y0.n460 0.00156143
R8566 Y0.n704 Y0.n703 0.00156143
R8567 Y0.n1059 Y0.n164 0.00156143
R8568 Y0.n1165 Y0.n113 0.00156143
R8569 Y0.n793 Y0.n792 0.00156143
R8570 Y0.n870 Y0.n869 0.00156143
R8571 Y0.n555 Y0.n554 0.00154762
R8572 Y0.n607 Y0.n606 0.00154762
R8573 Y0.n525 Y0.n402 0.00153931
R8574 Y0.n638 Y0.n361 0.00153931
R8575 Y0.n557 Y0.n556 0.00149509
R8576 Y0.n1170 Y0.n1169 0.00149509
R8577 Y0.n610 Y0.n370 0.00147297
R8578 Y0.n673 Y0.n347 0.00147297
R8579 Y0.n458 Y0.n426 0.00146905
R8580 Y0.n706 Y0.n705 0.00146905
R8581 Y0.n488 Y0.n413 0.00145086
R8582 Y0.n1214 Y0.n1213 0.00140663
R8583 Y0.n1335 Y0.n22 0.00140663
R8584 Y0.n493 Y0.n413 0.00140663
R8585 Y0.n674 Y0.n673 0.00140663
R8586 Y0.n589 Y0.n588 0.00139048
R8587 Y0.n556 Y0.n390 0.00138452
R8588 Y0.n605 Y0.n370 0.00138452
R8589 Y0.n450 Y0.n449 0.00136429
R8590 Y0.n566 Y0.n387 0.00136429
R8591 Y0.n572 Y0.n382 0.00136429
R8592 Y0.n526 Y0.n525 0.00134029
R8593 Y0.n643 Y0.n361 0.00134029
R8594 Y0.n598 Y0.n597 0.00133809
R8595 Y0.n715 Y0.n714 0.00133809
R8596 Y0.n460 Y0.n459 0.00131818
R8597 Y0.n704 Y0.n336 0.00131818
R8598 Y0.n1059 Y0.n1058 0.00131818
R8599 Y0.n755 Y0.n316 0.00129607
R8600 Y0.n777 Y0.n311 0.00129607
R8601 Y0.n832 Y0.n831 0.00129607
R8602 Y0.n855 Y0.n292 0.00129607
R8603 Y0.n473 Y0.n472 0.00128571
R8604 Y0.n691 Y0.n342 0.00128571
R8605 Y0.n1239 Y0.n68 0.00125184
R8606 Y0.n1309 Y0.n1308 0.00125184
R8607 Y0.n526 Y0.n404 0.00125184
R8608 Y0.n587 Y0.n377 0.00125184
R8609 Y0.n643 Y0.n642 0.00125184
R8610 Y0.n451 Y0.n429 0.00122973
R8611 Y0.n568 Y0.n567 0.00122973
R8612 Y0.n386 Y0.n383 0.00122973
R8613 Y0.n596 Y0.n374 0.00120762
R8614 Y0.n713 Y0.n333 0.00120762
R8615 Y0.n546 Y0.n395 0.00120714
R8616 Y0.n623 Y0.n366 0.00120714
R8617 Y0.n493 Y0.n492 0.0011855
R8618 Y0.n674 Y0.n349 0.0011855
R8619 Y0.n471 Y0.n420 0.00116339
R8620 Y0.n693 Y0.n692 0.00116339
R8621 Y0.n989 Y0.n198 0.00114865
R8622 Y0.n1100 Y0.n145 0.00114865
R8623 Y0.n745 Y0.n744 0.00114865
R8624 Y0.n819 Y0.n271 0.00114865
R8625 Y0.n663 Y0.n352 0.00112857
R8626 Y0.n610 Y0.n609 0.00111916
R8627 Y0.n506 Y0.n409 0.00110238
R8628 Y0.n1232 Y0.n1231 0.00109705
R8629 Y0.n38 Y0.n32 0.00109705
R8630 Y0.n545 Y0.n396 0.00109705
R8631 Y0.n557 Y0.n392 0.00109705
R8632 Y0.n622 Y0.n621 0.00109705
R8633 Y0.n1170 Y0.n112 0.00109705
R8634 Y0.n773 Y0.n772 0.00105283
R8635 Y0.n851 Y0.n850 0.00105283
R8636 Y0.n1358 Y0.n16 0.00105283
R8637 Y0.n1270 Y0.n53 0.00104054
R8638 Y0.n576 Y0.n226 0.00104054
R8639 Y0.n462 Y0.n461 0.00103071
R8640 Y0.n662 Y0.n353 0.00103071
R8641 Y0.n703 Y0.n338 0.00103071
R8642 Y0.n439 Y0.n432 0.00103071
R8643 Y0.n974 Y0.n973 0.00103071
R8644 Y0.n1085 Y0.n1084 0.00103071
R8645 Y0.n718 Y0.n331 0.00103071
R8646 Y0.n758 Y0.n757 0.00103071
R8647 Y0.n838 Y0.n837 0.00103071
R8648 Y0.n505 Y0.n504 0.0010086
R8649 Y0.n578 Y0.n577 0.000964373
R8650 Y0.n586 Y0.n379 0.000964373
R8651 Y0.n434 Y0.n433 0.000964373
R8652 Y0.n105 Y0.n102 0.000964373
R8653 Y0.n725 Y0.n328 0.000964373
R8654 Y0.n81 Y0.n78 0.00094226
R8655 Y0.n1315 Y0.n24 0.00094226
R8656 Y0.n199 Y0.n194 0.000932432
R8657 Y0.n146 Y0.n141 0.000932432
R8658 Y0.n749 Y0.n251 0.000932432
R8659 Y0.n825 Y0.n272 0.000932432
R8660 Y0.n444 Y0.n431 0.000898034
R8661 Y0.n695 Y0.n694 0.000898034
R8662 Y0.n470 Y0.n422 0.000875921
R8663 Y0.n728 Y0.n330 0.000853808
R8664 Y0.n1157 Y0.n1156 0.000831695
R8665 Y0.n1160 Y0.n1159 0.000814286
R8666 Y0.n544 Y0.n394 0.000809582
R8667 Y0.n620 Y0.n617 0.000809582
R8668 Y0.n1246 Y0.n1245 0.000787469
R8669 Y0.n1284 Y0.n1283 0.000787469
R8670 Y0.n1000 Y0.n999 0.000787469
R8671 Y0.n1111 Y0.n1110 0.000787469
R8672 Y0.n1158 Y0.n114 0.000765356
R8673 Y0.n743 Y0.n318 0.000765356
R8674 Y0.n788 Y0.n308 0.000765356
R8675 Y0.n821 Y0.n820 0.000765356
R8676 Y0.n865 Y0.n285 0.000765356
R8677 Y0.n661 Y0.n351 0.000743243
R8678 Y0.n503 Y0.n500 0.00072113
R8679 Y0.n95 Y0.n94 0.000716216
R8680 Y0.n1345 Y0.n19 0.000716216
R8681 Y0.n469 Y0.n212 0.000716216
R8682 Y0.n339 Y0.n241 0.000716216
R8683 Y0.n514 Y0.n406 0.000676904
R8684 Y0.n1199 Y0.n1198 0.000654791
R8685 Y0.n1343 Y0.n18 0.000654791
R8686 Y0.n651 Y0.n650 0.000654791
R8687 Y0.n631 Y0.n363 0.000588452
R8688 Y0.n534 Y0.n533 0.000566339
R8689 Y0.n1189 Y0.n101 0.000522113
R8690 Y0.n484 Y0.n483 0.000522113
R8691 Y1.n1377 Y1 18.2264
R8692 Y1.n1376 Y1.n1373 15.1827
R8693 Y1.n1375 Y1.n1374 15.0005
R8694 Y1 Y1.n1376 9.43874
R8695 Y1.n1377 Y1 9.19322
R8696 Y1.n1351 Y1.n19 2.2505
R8697 Y1.n34 Y1.n16 2.2505
R8698 Y1.n1357 Y1.n14 2.2505
R8699 Y1.n1303 Y1.n11 2.2505
R8700 Y1.n1363 Y1.n9 2.2505
R8701 Y1.n1283 Y1.n6 2.2505
R8702 Y1.n1369 Y1.n4 2.2505
R8703 Y1.n1370 Y1.n3 2.2505
R8704 Y1.n1254 Y1.n1253 2.2505
R8705 Y1.n1249 Y1.n1248 2.2505
R8706 Y1.n1227 Y1.n1226 2.2505
R8707 Y1.n1222 Y1.n1221 2.2505
R8708 Y1.n1208 Y1.n1207 2.2505
R8709 Y1.n1203 Y1.n1202 2.2505
R8710 Y1.n1183 Y1.n1182 2.2505
R8711 Y1.n950 Y1.n198 2.2505
R8712 Y1.n948 Y1.n200 2.2505
R8713 Y1.n944 Y1.n203 2.2505
R8714 Y1.n942 Y1.n205 2.2505
R8715 Y1.n938 Y1.n208 2.2505
R8716 Y1.n936 Y1.n210 2.2505
R8717 Y1.n932 Y1.n213 2.2505
R8718 Y1.n930 Y1.n215 2.2505
R8719 Y1.n361 Y1.n216 2.2505
R8720 Y1.n925 Y1.n219 2.2505
R8721 Y1.n617 Y1.n221 2.2505
R8722 Y1.n919 Y1.n224 2.2505
R8723 Y1.n664 Y1.n226 2.2505
R8724 Y1.n913 Y1.n229 2.2505
R8725 Y1.n320 Y1.n231 2.2505
R8726 Y1.n951 Y1.n950 2.2505
R8727 Y1.n948 Y1.n947 2.2505
R8728 Y1.n945 Y1.n944 2.2505
R8729 Y1.n942 Y1.n941 2.2505
R8730 Y1.n939 Y1.n938 2.2505
R8731 Y1.n936 Y1.n935 2.2505
R8732 Y1.n933 Y1.n932 2.2505
R8733 Y1.n930 Y1.n929 2.2505
R8734 Y1.n928 Y1.n216 2.2505
R8735 Y1.n925 Y1.n217 2.2505
R8736 Y1.n922 Y1.n221 2.2505
R8737 Y1.n919 Y1.n222 2.2505
R8738 Y1.n916 Y1.n226 2.2505
R8739 Y1.n913 Y1.n227 2.2505
R8740 Y1.n910 Y1.n231 2.2505
R8741 Y1.n1179 Y1.n1178 2.2505
R8742 Y1.n92 Y1.n91 2.2505
R8743 Y1.n1163 Y1.n1162 2.2505
R8744 Y1.n1161 Y1.n99 2.2505
R8745 Y1.n1160 Y1.n1159 2.2505
R8746 Y1.n101 Y1.n100 2.2505
R8747 Y1.n1116 Y1.n1115 2.2505
R8748 Y1.n1117 Y1.n1114 2.2505
R8749 Y1.n1118 Y1.n1113 2.2505
R8750 Y1.n1112 Y1.n116 2.2505
R8751 Y1.n1111 Y1.n1110 2.2505
R8752 Y1.n118 Y1.n117 2.2505
R8753 Y1.n1075 Y1.n1074 2.2505
R8754 Y1.n1082 Y1.n1073 2.2505
R8755 Y1.n1083 Y1.n1072 2.2505
R8756 Y1.n1071 Y1.n134 2.2505
R8757 Y1.n1070 Y1.n1069 2.2505
R8758 Y1.n136 Y1.n135 2.2505
R8759 Y1.n1053 Y1.n1052 2.2505
R8760 Y1.n1051 Y1.n151 2.2505
R8761 Y1.n1050 Y1.n1049 2.2505
R8762 Y1.n153 Y1.n152 2.2505
R8763 Y1.n1009 Y1.n1008 2.2505
R8764 Y1.n1016 Y1.n1007 2.2505
R8765 Y1.n1017 Y1.n1006 2.2505
R8766 Y1.n1005 Y1.n170 2.2505
R8767 Y1.n1004 Y1.n1003 2.2505
R8768 Y1.n172 Y1.n171 2.2505
R8769 Y1.n982 Y1.n981 2.2505
R8770 Y1.n980 Y1.n183 2.2505
R8771 Y1.n979 Y1.n978 2.2505
R8772 Y1.n185 Y1.n184 2.2505
R8773 Y1.n955 Y1.n954 2.2505
R8774 Y1.n956 Y1.n953 2.2505
R8775 Y1.n957 Y1.n956 2.2505
R8776 Y1.n955 Y1.n189 2.2505
R8777 Y1.n969 Y1.n185 2.2505
R8778 Y1.n978 Y1.n977 2.2505
R8779 Y1.n187 Y1.n183 2.2505
R8780 Y1.n983 Y1.n982 2.2505
R8781 Y1.n994 Y1.n172 2.2505
R8782 Y1.n1003 Y1.n1002 2.2505
R8783 Y1.n170 Y1.n167 2.2505
R8784 Y1.n1018 Y1.n1017 2.2505
R8785 Y1.n1016 Y1.n1015 2.2505
R8786 Y1.n1009 Y1.n158 2.2505
R8787 Y1.n1031 Y1.n153 2.2505
R8788 Y1.n1049 Y1.n1048 2.2505
R8789 Y1.n1037 Y1.n151 2.2505
R8790 Y1.n1054 Y1.n1053 2.2505
R8791 Y1.n1056 Y1.n136 2.2505
R8792 Y1.n1069 Y1.n1068 2.2505
R8793 Y1.n138 Y1.n134 2.2505
R8794 Y1.n1084 Y1.n1083 2.2505
R8795 Y1.n1082 Y1.n1081 2.2505
R8796 Y1.n1078 Y1.n1075 2.2505
R8797 Y1.n1095 Y1.n118 2.2505
R8798 Y1.n1110 Y1.n1109 2.2505
R8799 Y1.n1101 Y1.n116 2.2505
R8800 Y1.n1119 Y1.n1118 2.2505
R8801 Y1.n1117 Y1.n111 2.2505
R8802 Y1.n1116 Y1.n108 2.2505
R8803 Y1.n1135 Y1.n101 2.2505
R8804 Y1.n1159 Y1.n1158 2.2505
R8805 Y1.n1142 Y1.n99 2.2505
R8806 Y1.n1164 Y1.n1163 2.2505
R8807 Y1.n1166 Y1.n92 2.2505
R8808 Y1.n1178 Y1.n1177 2.2505
R8809 Y1.n907 Y1.n234 2.2505
R8810 Y1.n906 Y1.n235 2.2505
R8811 Y1.n905 Y1.n236 2.2505
R8812 Y1.n733 Y1.n237 2.2505
R8813 Y1.n901 Y1.n239 2.2505
R8814 Y1.n900 Y1.n240 2.2505
R8815 Y1.n899 Y1.n241 2.2505
R8816 Y1.n748 Y1.n242 2.2505
R8817 Y1.n895 Y1.n244 2.2505
R8818 Y1.n894 Y1.n245 2.2505
R8819 Y1.n893 Y1.n246 2.2505
R8820 Y1.n298 Y1.n247 2.2505
R8821 Y1.n889 Y1.n249 2.2505
R8822 Y1.n888 Y1.n250 2.2505
R8823 Y1.n887 Y1.n251 2.2505
R8824 Y1.n787 Y1.n252 2.2505
R8825 Y1.n883 Y1.n254 2.2505
R8826 Y1.n882 Y1.n255 2.2505
R8827 Y1.n881 Y1.n256 2.2505
R8828 Y1.n805 Y1.n257 2.2505
R8829 Y1.n877 Y1.n259 2.2505
R8830 Y1.n876 Y1.n260 2.2505
R8831 Y1.n875 Y1.n261 2.2505
R8832 Y1.n822 Y1.n262 2.2505
R8833 Y1.n871 Y1.n264 2.2505
R8834 Y1.n870 Y1.n265 2.2505
R8835 Y1.n869 Y1.n266 2.2505
R8836 Y1.n281 Y1.n267 2.2505
R8837 Y1.n865 Y1.n269 2.2505
R8838 Y1.n864 Y1.n270 2.2505
R8839 Y1.n863 Y1.n861 2.2505
R8840 Y1.n275 Y1.n23 2.2505
R8841 Y1.n1346 Y1.n1345 2.2505
R8842 Y1.n25 Y1.n20 2.2505
R8843 Y1.n1348 Y1.n20 2.2505
R8844 Y1.n1347 Y1.n1346 2.2505
R8845 Y1.n23 Y1.n22 2.2505
R8846 Y1.n863 Y1.n862 2.2505
R8847 Y1.n864 Y1.n268 2.2505
R8848 Y1.n866 Y1.n865 2.2505
R8849 Y1.n867 Y1.n267 2.2505
R8850 Y1.n869 Y1.n868 2.2505
R8851 Y1.n870 Y1.n263 2.2505
R8852 Y1.n872 Y1.n871 2.2505
R8853 Y1.n873 Y1.n262 2.2505
R8854 Y1.n875 Y1.n874 2.2505
R8855 Y1.n876 Y1.n258 2.2505
R8856 Y1.n878 Y1.n877 2.2505
R8857 Y1.n879 Y1.n257 2.2505
R8858 Y1.n881 Y1.n880 2.2505
R8859 Y1.n882 Y1.n253 2.2505
R8860 Y1.n884 Y1.n883 2.2505
R8861 Y1.n885 Y1.n252 2.2505
R8862 Y1.n887 Y1.n886 2.2505
R8863 Y1.n888 Y1.n248 2.2505
R8864 Y1.n890 Y1.n889 2.2505
R8865 Y1.n891 Y1.n247 2.2505
R8866 Y1.n893 Y1.n892 2.2505
R8867 Y1.n894 Y1.n243 2.2505
R8868 Y1.n896 Y1.n895 2.2505
R8869 Y1.n897 Y1.n242 2.2505
R8870 Y1.n899 Y1.n898 2.2505
R8871 Y1.n900 Y1.n238 2.2505
R8872 Y1.n902 Y1.n901 2.2505
R8873 Y1.n903 Y1.n237 2.2505
R8874 Y1.n905 Y1.n904 2.2505
R8875 Y1.n906 Y1.n233 2.2505
R8876 Y1.n908 Y1.n907 2.2505
R8877 Y1.n1351 Y1.n17 2.2505
R8878 Y1.n1354 Y1.n16 2.2505
R8879 Y1.n1357 Y1.n12 2.2505
R8880 Y1.n1360 Y1.n11 2.2505
R8881 Y1.n1363 Y1.n7 2.2505
R8882 Y1.n1366 Y1.n6 2.2505
R8883 Y1.n1369 Y1.n1 2.2505
R8884 Y1.n1371 Y1.n1370 2.2505
R8885 Y1.n1253 Y1.n1252 2.2505
R8886 Y1.n1250 Y1.n1249 2.2505
R8887 Y1.n1226 Y1.n1225 2.2505
R8888 Y1.n1223 Y1.n1222 2.2505
R8889 Y1.n1207 Y1.n1206 2.2505
R8890 Y1.n1204 Y1.n1203 2.2505
R8891 Y1.n1182 Y1.n1181 2.2505
R8892 Y1.n29 Y1.n28 2.2005
R8893 Y1.n1185 Y1.n1184 2.2005
R8894 Y1.n1186 Y1.n87 2.2005
R8895 Y1.n1189 Y1.n1188 2.2005
R8896 Y1.n1191 Y1.n86 2.2005
R8897 Y1.n1193 Y1.n1192 2.2005
R8898 Y1.n82 Y1.n79 2.2005
R8899 Y1.n1201 Y1.n1200 2.2005
R8900 Y1.n84 Y1.n81 2.2005
R8901 Y1.n83 Y1.n75 2.2005
R8902 Y1.n1210 Y1.n1209 2.2005
R8903 Y1.n1211 Y1.n73 2.2005
R8904 Y1.n1213 Y1.n1212 2.2005
R8905 Y1.n1216 Y1.n1215 2.2005
R8906 Y1.n1217 Y1.n70 2.2005
R8907 Y1.n1220 Y1.n1219 2.2005
R8908 Y1.n71 Y1.n64 2.2005
R8909 Y1.n1231 Y1.n1230 2.2005
R8910 Y1.n1229 Y1.n65 2.2005
R8911 Y1.n1228 Y1.n62 2.2005
R8912 Y1.n1237 Y1.n61 2.2005
R8913 Y1.n1239 Y1.n1238 2.2005
R8914 Y1.n1242 Y1.n1241 2.2005
R8915 Y1.n1243 Y1.n57 2.2005
R8916 Y1.n1247 Y1.n1246 2.2005
R8917 Y1.n1245 Y1.n59 2.2005
R8918 Y1.n52 Y1.n51 2.2005
R8919 Y1.n1256 Y1.n1255 2.2005
R8920 Y1.n53 Y1.n49 2.2005
R8921 Y1.n1264 Y1.n48 2.2005
R8922 Y1.n1266 Y1.n1265 2.2005
R8923 Y1.n1268 Y1.n47 2.2005
R8924 Y1.n1270 Y1.n1269 2.2005
R8925 Y1.n1272 Y1.n1271 2.2005
R8926 Y1.n1274 Y1.n1273 2.2005
R8927 Y1.n1276 Y1.n1275 2.2005
R8928 Y1.n1278 Y1.n1277 2.2005
R8929 Y1.n1279 Y1.n44 2.2005
R8930 Y1.n1282 Y1.n1281 2.2005
R8931 Y1.n1284 Y1.n43 2.2005
R8932 Y1.n1286 Y1.n1285 2.2005
R8933 Y1.n1289 Y1.n1288 2.2005
R8934 Y1.n1287 Y1.n41 2.2005
R8935 Y1.n1295 Y1.n1294 2.2005
R8936 Y1.n1296 Y1.n40 2.2005
R8937 Y1.n1298 Y1.n1297 2.2005
R8938 Y1.n1301 Y1.n1300 2.2005
R8939 Y1.n1302 Y1.n39 2.2005
R8940 Y1.n1306 Y1.n1305 2.2005
R8941 Y1.n1304 Y1.n37 2.2005
R8942 Y1.n1314 Y1.n1313 2.2005
R8943 Y1.n1316 Y1.n1315 2.2005
R8944 Y1.n1318 Y1.n1317 2.2005
R8945 Y1.n1320 Y1.n1319 2.2005
R8946 Y1.n1322 Y1.n1321 2.2005
R8947 Y1.n1324 Y1.n1323 2.2005
R8948 Y1.n1327 Y1.n1326 2.2005
R8949 Y1.n1328 Y1.n33 2.2005
R8950 Y1.n1330 Y1.n1329 2.2005
R8951 Y1.n1332 Y1.n1331 2.2005
R8952 Y1.n1334 Y1.n1333 2.2005
R8953 Y1.n712 Y1.n711 2.2005
R8954 Y1.n700 Y1.n699 2.2005
R8955 Y1.n698 Y1.n697 2.2005
R8956 Y1.n691 Y1.n690 2.2005
R8957 Y1.n689 Y1.n688 2.2005
R8958 Y1.n682 Y1.n327 2.2005
R8959 Y1.n673 Y1.n331 2.2005
R8960 Y1.n675 Y1.n674 2.2005
R8961 Y1.n665 Y1.n333 2.2005
R8962 Y1.n667 Y1.n666 2.2005
R8963 Y1.n663 Y1.n662 2.2005
R8964 Y1.n655 Y1.n336 2.2005
R8965 Y1.n649 Y1.n648 2.2005
R8966 Y1.n647 Y1.n646 2.2005
R8967 Y1.n642 Y1.n641 2.2005
R8968 Y1.n640 Y1.n639 2.2005
R8969 Y1.n634 Y1.n633 2.2005
R8970 Y1.n632 Y1.n631 2.2005
R8971 Y1.n625 Y1.n348 2.2005
R8972 Y1.n619 Y1.n618 2.2005
R8973 Y1.n616 Y1.n615 2.2005
R8974 Y1.n606 Y1.n353 2.2005
R8975 Y1.n608 Y1.n607 2.2005
R8976 Y1.n601 Y1.n600 2.2005
R8977 Y1.n599 Y1.n598 2.2005
R8978 Y1.n592 Y1.n591 2.2005
R8979 Y1.n590 Y1.n589 2.2005
R8980 Y1.n583 Y1.n582 2.2005
R8981 Y1.n581 Y1.n580 2.2005
R8982 Y1.n574 Y1.n573 2.2005
R8983 Y1.n572 Y1.n571 2.2005
R8984 Y1.n565 Y1.n564 2.2005
R8985 Y1.n563 Y1.n562 2.2005
R8986 Y1.n557 Y1.n372 2.2005
R8987 Y1.n548 Y1.n376 2.2005
R8988 Y1.n550 Y1.n549 2.2005
R8989 Y1.n546 Y1.n545 2.2005
R8990 Y1.n538 Y1.n379 2.2005
R8991 Y1.n532 Y1.n531 2.2005
R8992 Y1.n530 Y1.n529 2.2005
R8993 Y1.n525 Y1.n524 2.2005
R8994 Y1.n523 Y1.n522 2.2005
R8995 Y1.n517 Y1.n516 2.2005
R8996 Y1.n515 Y1.n514 2.2005
R8997 Y1.n508 Y1.n391 2.2005
R8998 Y1.n502 Y1.n501 2.2005
R8999 Y1.n499 Y1.n498 2.2005
R9000 Y1.n489 Y1.n396 2.2005
R9001 Y1.n491 Y1.n490 2.2005
R9002 Y1.n484 Y1.n483 2.2005
R9003 Y1.n482 Y1.n481 2.2005
R9004 Y1.n475 Y1.n474 2.2005
R9005 Y1.n473 Y1.n472 2.2005
R9006 Y1.n466 Y1.n465 2.2005
R9007 Y1.n464 Y1.n463 2.2005
R9008 Y1.n458 Y1.n457 2.2005
R9009 Y1.n456 Y1.n455 2.2005
R9010 Y1.n449 Y1.n411 2.2005
R9011 Y1.n440 Y1.n415 2.2005
R9012 Y1.n442 Y1.n441 2.2005
R9013 Y1.n435 Y1.n434 2.2005
R9014 Y1.n421 Y1.n195 2.2005
R9015 Y1.n958 Y1.n194 2.2005
R9016 Y1.n960 Y1.n959 2.2005
R9017 Y1.n967 Y1.n966 2.2005
R9018 Y1.n968 Y1.n188 2.2005
R9019 Y1.n971 Y1.n970 2.2005
R9020 Y1.n973 Y1.n186 2.2005
R9021 Y1.n976 Y1.n975 2.2005
R9022 Y1.n182 Y1.n181 2.2005
R9023 Y1.n986 Y1.n984 2.2005
R9024 Y1.n177 Y1.n176 2.2005
R9025 Y1.n993 Y1.n992 2.2005
R9026 Y1.n996 Y1.n995 2.2005
R9027 Y1.n998 Y1.n173 2.2005
R9028 Y1.n1001 Y1.n1000 2.2005
R9029 Y1.n174 Y1.n165 2.2005
R9030 Y1.n1021 Y1.n1020 2.2005
R9031 Y1.n1019 Y1.n166 2.2005
R9032 Y1.n169 Y1.n168 2.2005
R9033 Y1.n1011 Y1.n1010 2.2005
R9034 Y1.n1014 Y1.n1013 2.2005
R9035 Y1.n1012 Y1.n159 2.2005
R9036 Y1.n1029 Y1.n1028 2.2005
R9037 Y1.n1030 Y1.n157 2.2005
R9038 Y1.n1033 Y1.n1032 2.2005
R9039 Y1.n1035 Y1.n154 2.2005
R9040 Y1.n1047 Y1.n1046 2.2005
R9041 Y1.n1044 Y1.n155 2.2005
R9042 Y1.n1039 Y1.n1038 2.2005
R9043 Y1.n150 Y1.n148 2.2005
R9044 Y1.n1059 Y1.n1058 2.2005
R9045 Y1.n1057 Y1.n149 2.2005
R9046 Y1.n1055 Y1.n145 2.2005
R9047 Y1.n1064 Y1.n137 2.2005
R9048 Y1.n1067 Y1.n1066 2.2005
R9049 Y1.n140 Y1.n139 2.2005
R9050 Y1.n132 Y1.n130 2.2005
R9051 Y1.n1086 Y1.n1085 2.2005
R9052 Y1.n133 Y1.n131 2.2005
R9053 Y1.n1077 Y1.n1076 2.2005
R9054 Y1.n1080 Y1.n1079 2.2005
R9055 Y1.n125 Y1.n123 2.2005
R9056 Y1.n1094 Y1.n1093 2.2005
R9057 Y1.n1097 Y1.n1096 2.2005
R9058 Y1.n1099 Y1.n119 2.2005
R9059 Y1.n1108 Y1.n1107 2.2005
R9060 Y1.n1105 Y1.n120 2.2005
R9061 Y1.n1103 Y1.n1102 2.2005
R9062 Y1.n115 Y1.n114 2.2005
R9063 Y1.n1122 Y1.n1121 2.2005
R9064 Y1.n1120 Y1.n112 2.2005
R9065 Y1.n1128 Y1.n1127 2.2005
R9066 Y1.n1130 Y1.n1129 2.2005
R9067 Y1.n1133 Y1.n1132 2.2005
R9068 Y1.n1134 Y1.n107 2.2005
R9069 Y1.n1137 Y1.n1136 2.2005
R9070 Y1.n104 Y1.n102 2.2005
R9071 Y1.n1157 Y1.n1156 2.2005
R9072 Y1.n1140 Y1.n103 2.2005
R9073 Y1.n1144 Y1.n1143 2.2005
R9074 Y1.n1146 Y1.n98 2.2005
R9075 Y1.n1165 Y1.n97 2.2005
R9076 Y1.n1168 Y1.n1167 2.2005
R9077 Y1.n94 Y1.n93 2.2005
R9078 Y1.n1176 Y1.n1175 2.2005
R9079 Y1.n714 Y1.n713 2.2005
R9080 Y1.n723 Y1.n722 2.2005
R9081 Y1.n725 Y1.n724 2.2005
R9082 Y1.n727 Y1.n726 2.2005
R9083 Y1.n729 Y1.n728 2.2005
R9084 Y1.n730 Y1.n307 2.2005
R9085 Y1.n732 Y1.n731 2.2005
R9086 Y1.n735 Y1.n734 2.2005
R9087 Y1.n737 Y1.n736 2.2005
R9088 Y1.n739 Y1.n738 2.2005
R9089 Y1.n741 Y1.n740 2.2005
R9090 Y1.n743 Y1.n742 2.2005
R9091 Y1.n744 Y1.n303 2.2005
R9092 Y1.n747 Y1.n746 2.2005
R9093 Y1.n749 Y1.n302 2.2005
R9094 Y1.n751 Y1.n750 2.2005
R9095 Y1.n754 Y1.n753 2.2005
R9096 Y1.n752 Y1.n300 2.2005
R9097 Y1.n762 Y1.n761 2.2005
R9098 Y1.n764 Y1.n763 2.2005
R9099 Y1.n766 Y1.n765 2.2005
R9100 Y1.n768 Y1.n767 2.2005
R9101 Y1.n770 Y1.n769 2.2005
R9102 Y1.n772 Y1.n771 2.2005
R9103 Y1.n774 Y1.n773 2.2005
R9104 Y1.n776 Y1.n775 2.2005
R9105 Y1.n778 Y1.n777 2.2005
R9106 Y1.n780 Y1.n779 2.2005
R9107 Y1.n294 Y1.n293 2.2005
R9108 Y1.n786 Y1.n785 2.2005
R9109 Y1.n788 Y1.n292 2.2005
R9110 Y1.n790 Y1.n789 2.2005
R9111 Y1.n792 Y1.n791 2.2005
R9112 Y1.n794 Y1.n793 2.2005
R9113 Y1.n796 Y1.n795 2.2005
R9114 Y1.n798 Y1.n797 2.2005
R9115 Y1.n290 Y1.n289 2.2005
R9116 Y1.n804 Y1.n803 2.2005
R9117 Y1.n806 Y1.n288 2.2005
R9118 Y1.n808 Y1.n807 2.2005
R9119 Y1.n811 Y1.n810 2.2005
R9120 Y1.n813 Y1.n812 2.2005
R9121 Y1.n815 Y1.n814 2.2005
R9122 Y1.n286 Y1.n285 2.2005
R9123 Y1.n821 Y1.n820 2.2005
R9124 Y1.n823 Y1.n284 2.2005
R9125 Y1.n825 Y1.n824 2.2005
R9126 Y1.n828 Y1.n827 2.2005
R9127 Y1.n830 Y1.n829 2.2005
R9128 Y1.n833 Y1.n832 2.2005
R9129 Y1.n831 Y1.n282 2.2005
R9130 Y1.n840 Y1.n839 2.2005
R9131 Y1.n842 Y1.n841 2.2005
R9132 Y1.n844 Y1.n843 2.2005
R9133 Y1.n846 Y1.n845 2.2005
R9134 Y1.n848 Y1.n847 2.2005
R9135 Y1.n850 Y1.n849 2.2005
R9136 Y1.n852 Y1.n851 2.2005
R9137 Y1.n273 Y1.n271 2.2005
R9138 Y1.n860 Y1.n859 2.2005
R9139 Y1.n858 Y1.n272 2.2005
R9140 Y1.n277 Y1.n276 2.2005
R9141 Y1.n274 Y1.n24 2.2005
R9142 Y1.n1344 Y1.n1343 2.2005
R9143 Y1.n1342 Y1.n26 2.2005
R9144 Y1.n1352 Y1.n18 1.8005
R9145 Y1.n1356 Y1.n15 1.8005
R9146 Y1.n1358 Y1.n13 1.8005
R9147 Y1.n1362 Y1.n10 1.8005
R9148 Y1.n1364 Y1.n8 1.8005
R9149 Y1.n1368 Y1.n5 1.8005
R9150 Y1.n1267 Y1.n2 1.8005
R9151 Y1.n58 Y1.n54 1.8005
R9152 Y1.n1240 Y1.n56 1.8005
R9153 Y1.n67 Y1.n66 1.8005
R9154 Y1.n1214 Y1.n69 1.8005
R9155 Y1.n80 Y1.n76 1.8005
R9156 Y1.n1190 Y1.n78 1.8005
R9157 Y1.n949 Y1.n199 1.8005
R9158 Y1.n404 Y1.n201 1.8005
R9159 Y1.n943 Y1.n204 1.8005
R9160 Y1.n500 Y1.n206 1.8005
R9161 Y1.n937 Y1.n209 1.8005
R9162 Y1.n547 Y1.n211 1.8005
R9163 Y1.n931 Y1.n214 1.8005
R9164 Y1.n926 Y1.n218 1.8005
R9165 Y1.n924 Y1.n220 1.8005
R9166 Y1.n920 Y1.n223 1.8005
R9167 Y1.n918 Y1.n225 1.8005
R9168 Y1.n914 Y1.n228 1.8005
R9169 Y1.n912 Y1.n230 1.8005
R9170 Y1.n949 Y1.n197 1.8005
R9171 Y1.n946 Y1.n201 1.8005
R9172 Y1.n943 Y1.n202 1.8005
R9173 Y1.n940 Y1.n206 1.8005
R9174 Y1.n937 Y1.n207 1.8005
R9175 Y1.n934 Y1.n211 1.8005
R9176 Y1.n931 Y1.n212 1.8005
R9177 Y1.n927 Y1.n926 1.8005
R9178 Y1.n924 Y1.n923 1.8005
R9179 Y1.n921 Y1.n920 1.8005
R9180 Y1.n918 Y1.n917 1.8005
R9181 Y1.n915 Y1.n914 1.8005
R9182 Y1.n912 Y1.n911 1.8005
R9183 Y1.n1180 Y1.n90 1.8005
R9184 Y1.n90 Y1.n89 1.8005
R9185 Y1.n1350 Y1.n21 1.8005
R9186 Y1.n1350 Y1.n1349 1.8005
R9187 Y1.n1353 Y1.n1352 1.8005
R9188 Y1.n1356 Y1.n1355 1.8005
R9189 Y1.n1359 Y1.n1358 1.8005
R9190 Y1.n1362 Y1.n1361 1.8005
R9191 Y1.n1365 Y1.n1364 1.8005
R9192 Y1.n1368 Y1.n1367 1.8005
R9193 Y1.n2 Y1.n0 1.8005
R9194 Y1.n1251 Y1.n54 1.8005
R9195 Y1.n56 Y1.n55 1.8005
R9196 Y1.n1224 Y1.n67 1.8005
R9197 Y1.n69 Y1.n68 1.8005
R9198 Y1.n1205 Y1.n76 1.8005
R9199 Y1.n78 Y1.n77 1.8005
R9200 Y1.n952 Y1.n196 1.5005
R9201 Y1.n433 Y1.n196 1.5005
R9202 Y1.n715 Y1.n232 1.5005
R9203 Y1.n909 Y1.n232 1.5005
R9204 Y1.n719 Y1.n315 1.1125
R9205 Y1.n1150 Y1.n1145 1.10836
R9206 Y1.n1151 Y1.n1141 1.10443
R9207 Y1.n1174 Y1.n1173 1.10381
R9208 Y1.n718 Y1.n316 1.10372
R9209 Y1.n1155 Y1.n1154 1.10339
R9210 Y1.n97 Y1.n96 1.10272
R9211 Y1.n1149 Y1.n1146 1.10272
R9212 Y1.n1152 Y1.n1140 1.10272
R9213 Y1.n722 Y1.n721 1.10263
R9214 Y1.n725 Y1.n314 1.10263
R9215 Y1.n1336 Y1.n1335 1.1005
R9216 Y1.n1187 Y1.n85 1.1005
R9217 Y1.n1195 Y1.n1194 1.1005
R9218 Y1.n1199 Y1.n1198 1.1005
R9219 Y1.n1197 Y1.n74 1.1005
R9220 Y1.n1196 Y1.n72 1.1005
R9221 Y1.n1218 Y1.n63 1.1005
R9222 Y1.n1233 Y1.n1232 1.1005
R9223 Y1.n1236 Y1.n1235 1.1005
R9224 Y1.n1234 Y1.n60 1.1005
R9225 Y1.n1244 Y1.n50 1.1005
R9226 Y1.n1258 Y1.n1257 1.1005
R9227 Y1.n1263 Y1.n1262 1.1005
R9228 Y1.n1261 Y1.n47 1.1005
R9229 Y1.n1260 Y1.n46 1.1005
R9230 Y1.n1259 Y1.n45 1.1005
R9231 Y1.n1280 Y1.n42 1.1005
R9232 Y1.n1291 Y1.n1290 1.1005
R9233 Y1.n1293 Y1.n1292 1.1005
R9234 Y1.n1299 Y1.n38 1.1005
R9235 Y1.n1308 Y1.n1307 1.1005
R9236 Y1.n1312 Y1.n1311 1.1005
R9237 Y1.n1310 Y1.n36 1.1005
R9238 Y1.n1309 Y1.n35 1.1005
R9239 Y1.n1325 Y1.n32 1.1005
R9240 Y1.n1171 Y1.n88 1.1005
R9241 Y1.n961 Y1.n192 1.1005
R9242 Y1.n987 Y1.n179 1.1005
R9243 Y1.n1042 Y1.n1041 1.1005
R9244 Y1.n143 Y1.n142 1.1005
R9245 Y1.n1092 Y1.n1091 1.1005
R9246 Y1.n1170 Y1.n1169 1.1005
R9247 Y1.n1148 Y1.n1147 1.1005
R9248 Y1.n1153 Y1.n105 1.1005
R9249 Y1.n1139 Y1.n1138 1.1005
R9250 Y1.n1124 Y1.n1123 1.1005
R9251 Y1.n1090 Y1.n124 1.1005
R9252 Y1.n1088 Y1.n1087 1.1005
R9253 Y1.n144 Y1.n129 1.1005
R9254 Y1.n1061 Y1.n1060 1.1005
R9255 Y1.n1043 Y1.n147 1.1005
R9256 Y1.n1027 Y1.n1026 1.1005
R9257 Y1.n1023 Y1.n1022 1.1005
R9258 Y1.n989 Y1.n988 1.1005
R9259 Y1.n965 Y1.n964 1.1005
R9260 Y1.n963 Y1.n962 1.1005
R9261 Y1.n430 Y1.n423 1.1005
R9262 Y1.n429 Y1.n420 1.1005
R9263 Y1.n422 Y1.n193 1.1005
R9264 Y1.n432 Y1.n431 1.1005
R9265 Y1.n711 Y1.n710 1.1005
R9266 Y1.n702 Y1.n701 1.1005
R9267 Y1.n700 Y1.n322 1.1005
R9268 Y1.n697 Y1.n696 1.1005
R9269 Y1.n693 Y1.n692 1.1005
R9270 Y1.n686 Y1.n329 1.1005
R9271 Y1.n688 Y1.n687 1.1005
R9272 Y1.n685 Y1.n328 1.1005
R9273 Y1.n680 Y1.n679 1.1005
R9274 Y1.n669 Y1.n668 1.1005
R9275 Y1.n667 Y1.n334 1.1005
R9276 Y1.n659 Y1.n335 1.1005
R9277 Y1.n657 Y1.n656 1.1005
R9278 Y1.n655 Y1.n338 1.1005
R9279 Y1.n654 Y1.n653 1.1005
R9280 Y1.n341 Y1.n340 1.1005
R9281 Y1.n636 Y1.n345 1.1005
R9282 Y1.n635 Y1.n634 1.1005
R9283 Y1.n347 Y1.n346 1.1005
R9284 Y1.n627 Y1.n626 1.1005
R9285 Y1.n625 Y1.n350 1.1005
R9286 Y1.n624 Y1.n623 1.1005
R9287 Y1.n621 Y1.n620 1.1005
R9288 Y1.n615 Y1.n352 1.1005
R9289 Y1.n612 Y1.n353 1.1005
R9290 Y1.n609 Y1.n354 1.1005
R9291 Y1.n603 Y1.n355 1.1005
R9292 Y1.n602 Y1.n601 1.1005
R9293 Y1.n357 Y1.n356 1.1005
R9294 Y1.n594 Y1.n593 1.1005
R9295 Y1.n585 Y1.n584 1.1005
R9296 Y1.n583 Y1.n363 1.1005
R9297 Y1.n580 Y1.n579 1.1005
R9298 Y1.n576 Y1.n575 1.1005
R9299 Y1.n569 Y1.n369 1.1005
R9300 Y1.n571 Y1.n570 1.1005
R9301 Y1.n568 Y1.n368 1.1005
R9302 Y1.n560 Y1.n374 1.1005
R9303 Y1.n555 Y1.n554 1.1005
R9304 Y1.n553 Y1.n376 1.1005
R9305 Y1.n550 Y1.n377 1.1005
R9306 Y1.n544 Y1.n543 1.1005
R9307 Y1.n540 Y1.n539 1.1005
R9308 Y1.n538 Y1.n381 1.1005
R9309 Y1.n537 Y1.n536 1.1005
R9310 Y1.n384 Y1.n383 1.1005
R9311 Y1.n519 Y1.n388 1.1005
R9312 Y1.n518 Y1.n517 1.1005
R9313 Y1.n390 Y1.n389 1.1005
R9314 Y1.n510 Y1.n509 1.1005
R9315 Y1.n508 Y1.n393 1.1005
R9316 Y1.n507 Y1.n506 1.1005
R9317 Y1.n504 Y1.n503 1.1005
R9318 Y1.n498 Y1.n395 1.1005
R9319 Y1.n495 Y1.n396 1.1005
R9320 Y1.n492 Y1.n397 1.1005
R9321 Y1.n486 Y1.n398 1.1005
R9322 Y1.n485 Y1.n484 1.1005
R9323 Y1.n400 Y1.n399 1.1005
R9324 Y1.n477 Y1.n476 1.1005
R9325 Y1.n475 Y1.n402 1.1005
R9326 Y1.n469 Y1.n403 1.1005
R9327 Y1.n468 Y1.n405 1.1005
R9328 Y1.n467 Y1.n466 1.1005
R9329 Y1.n463 Y1.n462 1.1005
R9330 Y1.n460 Y1.n459 1.1005
R9331 Y1.n453 Y1.n413 1.1005
R9332 Y1.n455 Y1.n454 1.1005
R9333 Y1.n452 Y1.n412 1.1005
R9334 Y1.n447 Y1.n446 1.1005
R9335 Y1.n437 Y1.n417 1.1005
R9336 Y1.n436 Y1.n435 1.1005
R9337 Y1.n427 Y1.n426 1.1005
R9338 Y1.n428 Y1.n427 1.1005
R9339 Y1.n425 Y1.n420 1.1005
R9340 Y1.n419 Y1.n418 1.1005
R9341 Y1.n445 Y1.n415 1.1005
R9342 Y1.n444 Y1.n443 1.1005
R9343 Y1.n442 Y1.n416 1.1005
R9344 Y1.n439 Y1.n438 1.1005
R9345 Y1.n448 Y1.n414 1.1005
R9346 Y1.n451 Y1.n450 1.1005
R9347 Y1.n410 Y1.n409 1.1005
R9348 Y1.n461 Y1.n408 1.1005
R9349 Y1.n407 Y1.n406 1.1005
R9350 Y1.n471 Y1.n470 1.1005
R9351 Y1.n478 Y1.n401 1.1005
R9352 Y1.n480 Y1.n479 1.1005
R9353 Y1.n488 Y1.n487 1.1005
R9354 Y1.n494 Y1.n493 1.1005
R9355 Y1.n497 Y1.n496 1.1005
R9356 Y1.n505 Y1.n394 1.1005
R9357 Y1.n511 Y1.n392 1.1005
R9358 Y1.n513 Y1.n512 1.1005
R9359 Y1.n521 Y1.n520 1.1005
R9360 Y1.n529 Y1.n528 1.1005
R9361 Y1.n527 Y1.n385 1.1005
R9362 Y1.n526 Y1.n525 1.1005
R9363 Y1.n387 Y1.n386 1.1005
R9364 Y1.n534 Y1.n533 1.1005
R9365 Y1.n535 Y1.n382 1.1005
R9366 Y1.n541 Y1.n380 1.1005
R9367 Y1.n542 Y1.n378 1.1005
R9368 Y1.n552 Y1.n551 1.1005
R9369 Y1.n562 Y1.n561 1.1005
R9370 Y1.n559 Y1.n373 1.1005
R9371 Y1.n558 Y1.n557 1.1005
R9372 Y1.n556 Y1.n375 1.1005
R9373 Y1.n371 Y1.n370 1.1005
R9374 Y1.n567 Y1.n566 1.1005
R9375 Y1.n367 Y1.n366 1.1005
R9376 Y1.n577 Y1.n365 1.1005
R9377 Y1.n578 Y1.n364 1.1005
R9378 Y1.n592 Y1.n359 1.1005
R9379 Y1.n587 Y1.n360 1.1005
R9380 Y1.n589 Y1.n588 1.1005
R9381 Y1.n586 Y1.n362 1.1005
R9382 Y1.n595 Y1.n358 1.1005
R9383 Y1.n597 Y1.n596 1.1005
R9384 Y1.n605 Y1.n604 1.1005
R9385 Y1.n611 Y1.n610 1.1005
R9386 Y1.n614 Y1.n613 1.1005
R9387 Y1.n622 Y1.n351 1.1005
R9388 Y1.n628 Y1.n349 1.1005
R9389 Y1.n630 Y1.n629 1.1005
R9390 Y1.n638 Y1.n637 1.1005
R9391 Y1.n646 Y1.n645 1.1005
R9392 Y1.n644 Y1.n342 1.1005
R9393 Y1.n643 Y1.n642 1.1005
R9394 Y1.n344 Y1.n343 1.1005
R9395 Y1.n651 Y1.n650 1.1005
R9396 Y1.n652 Y1.n339 1.1005
R9397 Y1.n658 Y1.n337 1.1005
R9398 Y1.n661 Y1.n660 1.1005
R9399 Y1.n670 Y1.n333 1.1005
R9400 Y1.n678 Y1.n331 1.1005
R9401 Y1.n677 Y1.n676 1.1005
R9402 Y1.n675 Y1.n332 1.1005
R9403 Y1.n672 Y1.n671 1.1005
R9404 Y1.n681 Y1.n330 1.1005
R9405 Y1.n684 Y1.n683 1.1005
R9406 Y1.n326 Y1.n325 1.1005
R9407 Y1.n694 Y1.n324 1.1005
R9408 Y1.n695 Y1.n323 1.1005
R9409 Y1.n703 Y1.n321 1.1005
R9410 Y1.n709 Y1.n318 1.1005
R9411 Y1.n319 Y1.n317 1.1005
R9412 Y1.n706 Y1.n705 1.1005
R9413 Y1.n1340 Y1.n1339 1.1005
R9414 Y1.n1338 Y1.n31 1.1005
R9415 Y1.n1337 Y1.n31 1.1005
R9416 Y1.n708 Y1.n319 1.1005
R9417 Y1.n707 Y1.n706 1.1005
R9418 Y1.n1341 Y1.n30 1.1005
R9419 Y1.n855 Y1.n27 1.1005
R9420 Y1.n857 Y1.n856 1.1005
R9421 Y1.n854 Y1.n853 1.1005
R9422 Y1.n279 Y1.n278 1.1005
R9423 Y1.n836 Y1.n280 1.1005
R9424 Y1.n838 Y1.n837 1.1005
R9425 Y1.n835 Y1.n834 1.1005
R9426 Y1.n826 Y1.n283 1.1005
R9427 Y1.n819 Y1.n818 1.1005
R9428 Y1.n817 Y1.n816 1.1005
R9429 Y1.n809 Y1.n287 1.1005
R9430 Y1.n802 Y1.n801 1.1005
R9431 Y1.n800 Y1.n799 1.1005
R9432 Y1.n791 Y1.n291 1.1005
R9433 Y1.n784 Y1.n783 1.1005
R9434 Y1.n782 Y1.n781 1.1005
R9435 Y1.n296 Y1.n295 1.1005
R9436 Y1.n757 Y1.n297 1.1005
R9437 Y1.n758 Y1.n299 1.1005
R9438 Y1.n760 Y1.n759 1.1005
R9439 Y1.n756 Y1.n755 1.1005
R9440 Y1.n745 Y1.n301 1.1005
R9441 Y1.n310 Y1.n304 1.1005
R9442 Y1.n311 Y1.n305 1.1005
R9443 Y1.n312 Y1.n306 1.1005
R9444 Y1.n313 Y1.n308 1.1005
R9445 Y1.n720 Y1.n309 1.1005
R9446 Y1.n717 Y1.n716 1.1005
R9447 Y1.n433 Y1.n432 0.733833
R9448 Y1.n95 Y1.n89 0.733833
R9449 Y1.n1341 Y1.n21 0.733833
R9450 Y1.n716 Y1.n715 0.733833
R9451 Y1.n1091 Y1.n122 0.573769
R9452 Y1.n985 Y1.n179 0.573769
R9453 Y1.n142 Y1.n141 0.573695
R9454 Y1.n192 Y1.n190 0.573695
R9455 Y1.n1041 Y1.n1040 0.573346
R9456 Y1.n424 Y1.n420 0.550549
R9457 Y1.n704 Y1.n319 0.550549
R9458 Y1.n1090 Y1.n126 0.39244
R9459 Y1.n989 Y1.n178 0.39244
R9460 Y1.n1065 Y1.n129 0.389994
R9461 Y1.n963 Y1.n191 0.389994
R9462 Y1.n1045 Y1.n147 0.387191
R9463 Y1.n1131 Y1.n106 0.384705
R9464 Y1.n1025 Y1.n160 0.384705
R9465 Y1.n1100 Y1.n121 0.384705
R9466 Y1.n990 Y1.n175 0.384705
R9467 Y1.n1125 Y1.n110 0.382331
R9468 Y1.n1024 Y1.n163 0.382331
R9469 Y1.n1106 Y1.n113 0.382034
R9470 Y1.n997 Y1.n164 0.382034
R9471 Y1.n1089 Y1.n127 0.379547
R9472 Y1.n1036 Y1.n156 0.379547
R9473 Y1.n972 Y1.n180 0.379547
R9474 Y1.n1063 Y1.n1062 0.376968
R9475 Y1.n1062 Y1.n146 0.376876
R9476 Y1.n1089 Y1.n128 0.375976
R9477 Y1.n974 Y1.n180 0.375976
R9478 Y1.n1034 Y1.n156 0.375884
R9479 Y1.n1104 Y1.n113 0.374982
R9480 Y1.n999 Y1.n164 0.374982
R9481 Y1.n1126 Y1.n1125 0.374889
R9482 Y1.n1024 Y1.n162 0.374889
R9483 Y1.n109 Y1.n106 0.373984
R9484 Y1.n1025 Y1.n161 0.373984
R9485 Y1.n1098 Y1.n121 0.373891
R9486 Y1.n991 Y1.n990 0.373891
R9487 Y1 Y1.n1372 0.296734
R9488 Y1.n1172 Y1.n95 0.275034
R9489 Y1.n1376 Y1.n1375 0.189306
R9490 Y1.n1375 Y1 0.0513955
R9491 Y1.n1182 Y1.n78 0.0405
R9492 Y1.n1203 Y1.n78 0.0405
R9493 Y1.n1203 Y1.n76 0.0405
R9494 Y1.n1207 Y1.n76 0.0405
R9495 Y1.n1207 Y1.n69 0.0405
R9496 Y1.n1222 Y1.n69 0.0405
R9497 Y1.n1222 Y1.n67 0.0405
R9498 Y1.n1226 Y1.n67 0.0405
R9499 Y1.n1226 Y1.n56 0.0405
R9500 Y1.n1249 Y1.n56 0.0405
R9501 Y1.n1249 Y1.n54 0.0405
R9502 Y1.n1253 Y1.n54 0.0405
R9503 Y1.n1253 Y1.n2 0.0405
R9504 Y1.n1370 Y1.n2 0.0405
R9505 Y1.n1369 Y1.n1368 0.0405
R9506 Y1.n1368 Y1.n6 0.0405
R9507 Y1.n1364 Y1.n6 0.0405
R9508 Y1.n1364 Y1.n1363 0.0405
R9509 Y1.n1363 Y1.n1362 0.0405
R9510 Y1.n1362 Y1.n11 0.0405
R9511 Y1.n1358 Y1.n11 0.0405
R9512 Y1.n1358 Y1.n1357 0.0405
R9513 Y1.n1357 Y1.n1356 0.0405
R9514 Y1.n1356 Y1.n16 0.0405
R9515 Y1.n1352 Y1.n16 0.0405
R9516 Y1.n1352 Y1.n1351 0.0405
R9517 Y1.n950 Y1.n949 0.0405
R9518 Y1.n949 Y1.n948 0.0405
R9519 Y1.n948 Y1.n201 0.0405
R9520 Y1.n944 Y1.n201 0.0405
R9521 Y1.n944 Y1.n943 0.0405
R9522 Y1.n943 Y1.n942 0.0405
R9523 Y1.n942 Y1.n206 0.0405
R9524 Y1.n938 Y1.n206 0.0405
R9525 Y1.n938 Y1.n937 0.0405
R9526 Y1.n937 Y1.n936 0.0405
R9527 Y1.n936 Y1.n211 0.0405
R9528 Y1.n932 Y1.n211 0.0405
R9529 Y1.n932 Y1.n931 0.0405
R9530 Y1.n931 Y1.n930 0.0405
R9531 Y1.n926 Y1.n216 0.0405
R9532 Y1.n926 Y1.n925 0.0405
R9533 Y1.n925 Y1.n924 0.0405
R9534 Y1.n924 Y1.n221 0.0405
R9535 Y1.n920 Y1.n221 0.0405
R9536 Y1.n920 Y1.n919 0.0405
R9537 Y1.n919 Y1.n918 0.0405
R9538 Y1.n918 Y1.n226 0.0405
R9539 Y1.n914 Y1.n226 0.0405
R9540 Y1.n914 Y1.n913 0.0405
R9541 Y1.n913 Y1.n912 0.0405
R9542 Y1.n912 Y1.n231 0.0405
R9543 Y1.n951 Y1.n197 0.0405
R9544 Y1.n947 Y1.n197 0.0405
R9545 Y1.n947 Y1.n946 0.0405
R9546 Y1.n946 Y1.n945 0.0405
R9547 Y1.n945 Y1.n202 0.0405
R9548 Y1.n941 Y1.n202 0.0405
R9549 Y1.n941 Y1.n940 0.0405
R9550 Y1.n940 Y1.n939 0.0405
R9551 Y1.n939 Y1.n207 0.0405
R9552 Y1.n935 Y1.n207 0.0405
R9553 Y1.n935 Y1.n934 0.0405
R9554 Y1.n934 Y1.n933 0.0405
R9555 Y1.n933 Y1.n212 0.0405
R9556 Y1.n929 Y1.n212 0.0405
R9557 Y1.n928 Y1.n927 0.0405
R9558 Y1.n927 Y1.n217 0.0405
R9559 Y1.n923 Y1.n217 0.0405
R9560 Y1.n923 Y1.n922 0.0405
R9561 Y1.n922 Y1.n921 0.0405
R9562 Y1.n921 Y1.n222 0.0405
R9563 Y1.n917 Y1.n222 0.0405
R9564 Y1.n917 Y1.n916 0.0405
R9565 Y1.n916 Y1.n915 0.0405
R9566 Y1.n915 Y1.n227 0.0405
R9567 Y1.n911 Y1.n227 0.0405
R9568 Y1.n911 Y1.n910 0.0405
R9569 Y1.n1181 Y1.n77 0.0405
R9570 Y1.n1204 Y1.n77 0.0405
R9571 Y1.n1205 Y1.n1204 0.0405
R9572 Y1.n1206 Y1.n1205 0.0405
R9573 Y1.n1206 Y1.n68 0.0405
R9574 Y1.n1223 Y1.n68 0.0405
R9575 Y1.n1224 Y1.n1223 0.0405
R9576 Y1.n1225 Y1.n1224 0.0405
R9577 Y1.n1225 Y1.n55 0.0405
R9578 Y1.n1250 Y1.n55 0.0405
R9579 Y1.n1251 Y1.n1250 0.0405
R9580 Y1.n1252 Y1.n1251 0.0405
R9581 Y1.n1252 Y1.n0 0.0405
R9582 Y1.n1367 Y1.n1 0.0405
R9583 Y1.n1367 Y1.n1366 0.0405
R9584 Y1.n1366 Y1.n1365 0.0405
R9585 Y1.n1365 Y1.n7 0.0405
R9586 Y1.n1361 Y1.n7 0.0405
R9587 Y1.n1361 Y1.n1360 0.0405
R9588 Y1.n1360 Y1.n1359 0.0405
R9589 Y1.n1359 Y1.n12 0.0405
R9590 Y1.n1355 Y1.n12 0.0405
R9591 Y1.n1355 Y1.n1354 0.0405
R9592 Y1.n1354 Y1.n1353 0.0405
R9593 Y1.n1353 Y1.n17 0.0405
R9594 Y1.n1370 Y1.n1369 0.0360676
R9595 Y1.n930 Y1.n216 0.0360676
R9596 Y1.n929 Y1.n928 0.0360676
R9597 Y1.n954 Y1.n953 0.0360676
R9598 Y1.n954 Y1.n184 0.0360676
R9599 Y1.n979 Y1.n184 0.0360676
R9600 Y1.n980 Y1.n979 0.0360676
R9601 Y1.n981 Y1.n980 0.0360676
R9602 Y1.n981 Y1.n171 0.0360676
R9603 Y1.n1004 Y1.n171 0.0360676
R9604 Y1.n1005 Y1.n1004 0.0360676
R9605 Y1.n1006 Y1.n1005 0.0360676
R9606 Y1.n1007 Y1.n1006 0.0360676
R9607 Y1.n1008 Y1.n1007 0.0360676
R9608 Y1.n1008 Y1.n152 0.0360676
R9609 Y1.n1050 Y1.n152 0.0360676
R9610 Y1.n1051 Y1.n1050 0.0360676
R9611 Y1.n1052 Y1.n1051 0.0360676
R9612 Y1.n1052 Y1.n135 0.0360676
R9613 Y1.n1070 Y1.n135 0.0360676
R9614 Y1.n1071 Y1.n1070 0.0360676
R9615 Y1.n1072 Y1.n1071 0.0360676
R9616 Y1.n1073 Y1.n1072 0.0360676
R9617 Y1.n1074 Y1.n1073 0.0360676
R9618 Y1.n1074 Y1.n117 0.0360676
R9619 Y1.n1111 Y1.n117 0.0360676
R9620 Y1.n1112 Y1.n1111 0.0360676
R9621 Y1.n1113 Y1.n1112 0.0360676
R9622 Y1.n1114 Y1.n1113 0.0360676
R9623 Y1.n1115 Y1.n1114 0.0360676
R9624 Y1.n1115 Y1.n100 0.0360676
R9625 Y1.n1160 Y1.n100 0.0360676
R9626 Y1.n1161 Y1.n1160 0.0360676
R9627 Y1.n1162 Y1.n1161 0.0360676
R9628 Y1.n1162 Y1.n91 0.0360676
R9629 Y1.n1179 Y1.n91 0.0360676
R9630 Y1.n956 Y1.n955 0.0360676
R9631 Y1.n955 Y1.n185 0.0360676
R9632 Y1.n978 Y1.n185 0.0360676
R9633 Y1.n978 Y1.n183 0.0360676
R9634 Y1.n982 Y1.n183 0.0360676
R9635 Y1.n982 Y1.n172 0.0360676
R9636 Y1.n1003 Y1.n172 0.0360676
R9637 Y1.n1003 Y1.n170 0.0360676
R9638 Y1.n1017 Y1.n170 0.0360676
R9639 Y1.n1017 Y1.n1016 0.0360676
R9640 Y1.n1016 Y1.n1009 0.0360676
R9641 Y1.n1009 Y1.n153 0.0360676
R9642 Y1.n1049 Y1.n153 0.0360676
R9643 Y1.n1049 Y1.n151 0.0360676
R9644 Y1.n1053 Y1.n151 0.0360676
R9645 Y1.n1053 Y1.n136 0.0360676
R9646 Y1.n1069 Y1.n136 0.0360676
R9647 Y1.n1069 Y1.n134 0.0360676
R9648 Y1.n1083 Y1.n134 0.0360676
R9649 Y1.n1083 Y1.n1082 0.0360676
R9650 Y1.n1082 Y1.n1075 0.0360676
R9651 Y1.n1075 Y1.n118 0.0360676
R9652 Y1.n1110 Y1.n118 0.0360676
R9653 Y1.n1110 Y1.n116 0.0360676
R9654 Y1.n1118 Y1.n116 0.0360676
R9655 Y1.n1118 Y1.n1117 0.0360676
R9656 Y1.n1117 Y1.n1116 0.0360676
R9657 Y1.n1116 Y1.n101 0.0360676
R9658 Y1.n1159 Y1.n101 0.0360676
R9659 Y1.n1159 Y1.n99 0.0360676
R9660 Y1.n1163 Y1.n99 0.0360676
R9661 Y1.n1163 Y1.n92 0.0360676
R9662 Y1.n1178 Y1.n92 0.0360676
R9663 Y1.n907 Y1.n906 0.0360676
R9664 Y1.n906 Y1.n905 0.0360676
R9665 Y1.n905 Y1.n237 0.0360676
R9666 Y1.n901 Y1.n237 0.0360676
R9667 Y1.n901 Y1.n900 0.0360676
R9668 Y1.n900 Y1.n899 0.0360676
R9669 Y1.n899 Y1.n242 0.0360676
R9670 Y1.n895 Y1.n242 0.0360676
R9671 Y1.n895 Y1.n894 0.0360676
R9672 Y1.n894 Y1.n893 0.0360676
R9673 Y1.n893 Y1.n247 0.0360676
R9674 Y1.n889 Y1.n247 0.0360676
R9675 Y1.n889 Y1.n888 0.0360676
R9676 Y1.n888 Y1.n887 0.0360676
R9677 Y1.n887 Y1.n252 0.0360676
R9678 Y1.n883 Y1.n252 0.0360676
R9679 Y1.n883 Y1.n882 0.0360676
R9680 Y1.n882 Y1.n881 0.0360676
R9681 Y1.n881 Y1.n257 0.0360676
R9682 Y1.n877 Y1.n257 0.0360676
R9683 Y1.n877 Y1.n876 0.0360676
R9684 Y1.n876 Y1.n875 0.0360676
R9685 Y1.n875 Y1.n262 0.0360676
R9686 Y1.n871 Y1.n262 0.0360676
R9687 Y1.n871 Y1.n870 0.0360676
R9688 Y1.n870 Y1.n869 0.0360676
R9689 Y1.n869 Y1.n267 0.0360676
R9690 Y1.n865 Y1.n267 0.0360676
R9691 Y1.n865 Y1.n864 0.0360676
R9692 Y1.n864 Y1.n863 0.0360676
R9693 Y1.n863 Y1.n23 0.0360676
R9694 Y1.n1346 Y1.n23 0.0360676
R9695 Y1.n1346 Y1.n20 0.0360676
R9696 Y1.n908 Y1.n233 0.0360676
R9697 Y1.n904 Y1.n233 0.0360676
R9698 Y1.n904 Y1.n903 0.0360676
R9699 Y1.n903 Y1.n902 0.0360676
R9700 Y1.n902 Y1.n238 0.0360676
R9701 Y1.n898 Y1.n238 0.0360676
R9702 Y1.n898 Y1.n897 0.0360676
R9703 Y1.n897 Y1.n896 0.0360676
R9704 Y1.n896 Y1.n243 0.0360676
R9705 Y1.n892 Y1.n243 0.0360676
R9706 Y1.n892 Y1.n891 0.0360676
R9707 Y1.n891 Y1.n890 0.0360676
R9708 Y1.n890 Y1.n248 0.0360676
R9709 Y1.n886 Y1.n248 0.0360676
R9710 Y1.n886 Y1.n885 0.0360676
R9711 Y1.n885 Y1.n884 0.0360676
R9712 Y1.n884 Y1.n253 0.0360676
R9713 Y1.n880 Y1.n253 0.0360676
R9714 Y1.n880 Y1.n879 0.0360676
R9715 Y1.n879 Y1.n878 0.0360676
R9716 Y1.n878 Y1.n258 0.0360676
R9717 Y1.n874 Y1.n258 0.0360676
R9718 Y1.n874 Y1.n873 0.0360676
R9719 Y1.n873 Y1.n872 0.0360676
R9720 Y1.n872 Y1.n263 0.0360676
R9721 Y1.n868 Y1.n263 0.0360676
R9722 Y1.n868 Y1.n867 0.0360676
R9723 Y1.n867 Y1.n866 0.0360676
R9724 Y1.n866 Y1.n268 0.0360676
R9725 Y1.n862 Y1.n268 0.0360676
R9726 Y1.n862 Y1.n22 0.0360676
R9727 Y1.n1347 Y1.n22 0.0360676
R9728 Y1.n1348 Y1.n1347 0.0360676
R9729 Y1.n1371 Y1.n1 0.0360676
R9730 Y1.n1372 Y1.n1371 0.0248243
R9731 Y1 Y1.n1377 0.0245437
R9732 Y1.n1182 Y1.n90 0.0234189
R9733 Y1.n950 Y1.n196 0.0234189
R9734 Y1.n952 Y1.n951 0.0234189
R9735 Y1.n1181 Y1.n1180 0.0234189
R9736 Y1.n1351 Y1.n1350 0.0233108
R9737 Y1.n232 Y1.n231 0.0233108
R9738 Y1.n910 Y1.n909 0.0233108
R9739 Y1.n1349 Y1.n17 0.0233108
R9740 Y1.n953 Y1.n952 0.0227703
R9741 Y1.n956 Y1.n196 0.0227703
R9742 Y1.n907 Y1.n232 0.0227703
R9743 Y1.n909 Y1.n908 0.0227703
R9744 Y1.n1192 Y1.n79 0.0188784
R9745 Y1.n1201 Y1.n81 0.0188784
R9746 Y1.n1209 Y1.n75 0.0188784
R9747 Y1.n1213 Y1.n73 0.0188784
R9748 Y1.n1215 Y1.n70 0.0188784
R9749 Y1.n1229 Y1.n1228 0.0188784
R9750 Y1.n1239 Y1.n61 0.0188784
R9751 Y1.n1241 Y1.n57 0.0188784
R9752 Y1.n1247 Y1.n59 0.0188784
R9753 Y1.n1255 Y1.n52 0.0188784
R9754 Y1.n53 Y1.n48 0.0188784
R9755 Y1.n1269 Y1.n1268 0.0188784
R9756 Y1.n1273 Y1.n1272 0.0188784
R9757 Y1.n1277 Y1.n1276 0.0188784
R9758 Y1.n1282 Y1.n44 0.0188784
R9759 Y1.n1285 Y1.n1284 0.0188784
R9760 Y1.n1288 Y1.n1287 0.0188784
R9761 Y1.n1296 Y1.n1295 0.0188784
R9762 Y1.n1305 Y1.n1304 0.0188784
R9763 Y1.n1315 Y1.n1314 0.0188784
R9764 Y1.n1319 Y1.n1318 0.0188784
R9765 Y1.n1323 Y1.n1322 0.0188784
R9766 Y1.n1328 Y1.n1327 0.0188784
R9767 Y1.n457 Y1.n456 0.0188784
R9768 Y1.n465 Y1.n464 0.0188784
R9769 Y1.n474 Y1.n473 0.0188784
R9770 Y1.n483 Y1.n482 0.0188784
R9771 Y1.n490 Y1.n489 0.0188784
R9772 Y1.n516 Y1.n515 0.0188784
R9773 Y1.n524 Y1.n523 0.0188784
R9774 Y1.n531 Y1.n530 0.0188784
R9775 Y1.n546 Y1.n379 0.0188784
R9776 Y1.n549 Y1.n548 0.0188784
R9777 Y1.n563 Y1.n372 0.0188784
R9778 Y1.n573 Y1.n572 0.0188784
R9779 Y1.n582 Y1.n581 0.0188784
R9780 Y1.n591 Y1.n590 0.0188784
R9781 Y1.n600 Y1.n599 0.0188784
R9782 Y1.n607 Y1.n606 0.0188784
R9783 Y1.n618 Y1.n616 0.0188784
R9784 Y1.n632 Y1.n348 0.0188784
R9785 Y1.n648 Y1.n647 0.0188784
R9786 Y1.n663 Y1.n336 0.0188784
R9787 Y1.n666 Y1.n665 0.0188784
R9788 Y1.n674 Y1.n673 0.0188784
R9789 Y1.n689 Y1.n327 0.0188784
R9790 Y1.n433 Y1.n195 0.0188784
R9791 Y1.n959 Y1.n958 0.0188784
R9792 Y1.n968 Y1.n967 0.0188784
R9793 Y1.n970 Y1.n186 0.0188784
R9794 Y1.n1055 Y1.n137 0.0188784
R9795 Y1.n1067 Y1.n139 0.0188784
R9796 Y1.n1085 Y1.n132 0.0188784
R9797 Y1.n1077 Y1.n133 0.0188784
R9798 Y1.n715 Y1.n714 0.0188784
R9799 Y1.n724 Y1.n723 0.0188784
R9800 Y1.n728 Y1.n727 0.0188784
R9801 Y1.n732 Y1.n307 0.0188784
R9802 Y1.n793 Y1.n792 0.0188784
R9803 Y1.n797 Y1.n796 0.0188784
R9804 Y1.n804 Y1.n289 0.0188784
R9805 Y1.n807 Y1.n806 0.0188784
R9806 Y1.n1189 Y1.n87 0.0187703
R9807 Y1.n1192 Y1.n1191 0.0187703
R9808 Y1.n1220 Y1.n71 0.0187703
R9809 Y1.n1230 Y1.n1229 0.0187703
R9810 Y1.n1266 Y1.n48 0.0187703
R9811 Y1.n1297 Y1.n1296 0.0187703
R9812 Y1.n1302 Y1.n1301 0.0187703
R9813 Y1.n1329 Y1.n1328 0.0187703
R9814 Y1.n1333 Y1.n1332 0.0187703
R9815 Y1.n441 Y1.n440 0.0187703
R9816 Y1.n456 Y1.n411 0.0187703
R9817 Y1.n501 Y1.n499 0.0187703
R9818 Y1.n515 Y1.n391 0.0187703
R9819 Y1.n564 Y1.n563 0.0187703
R9820 Y1.n633 Y1.n632 0.0187703
R9821 Y1.n641 Y1.n640 0.0187703
R9822 Y1.n690 Y1.n689 0.0187703
R9823 Y1.n699 Y1.n698 0.0187703
R9824 Y1.n984 Y1.n182 0.0187703
R9825 Y1.n993 Y1.n176 0.0187703
R9826 Y1.n995 Y1.n173 0.0187703
R9827 Y1.n1001 Y1.n174 0.0187703
R9828 Y1.n1020 Y1.n1019 0.0187703
R9829 Y1.n1011 Y1.n169 0.0187703
R9830 Y1.n1014 Y1.n1012 0.0187703
R9831 Y1.n1030 Y1.n1029 0.0187703
R9832 Y1.n1032 Y1.n154 0.0187703
R9833 Y1.n1047 Y1.n155 0.0187703
R9834 Y1.n1038 Y1.n150 0.0187703
R9835 Y1.n1058 Y1.n1057 0.0187703
R9836 Y1.n1094 Y1.n123 0.0187703
R9837 Y1.n1096 Y1.n119 0.0187703
R9838 Y1.n1108 Y1.n120 0.0187703
R9839 Y1.n1102 Y1.n115 0.0187703
R9840 Y1.n1121 Y1.n1120 0.0187703
R9841 Y1.n1129 Y1.n1128 0.0187703
R9842 Y1.n1134 Y1.n1133 0.0187703
R9843 Y1.n1136 Y1.n102 0.0187703
R9844 Y1.n1157 Y1.n103 0.0187703
R9845 Y1.n1143 Y1.n98 0.0187703
R9846 Y1.n1167 Y1.n1165 0.0187703
R9847 Y1.n1176 Y1.n93 0.0187703
R9848 Y1.n738 Y1.n737 0.0187703
R9849 Y1.n742 Y1.n741 0.0187703
R9850 Y1.n747 Y1.n303 0.0187703
R9851 Y1.n750 Y1.n749 0.0187703
R9852 Y1.n753 Y1.n752 0.0187703
R9853 Y1.n763 Y1.n762 0.0187703
R9854 Y1.n767 Y1.n766 0.0187703
R9855 Y1.n771 Y1.n770 0.0187703
R9856 Y1.n775 Y1.n774 0.0187703
R9857 Y1.n779 Y1.n778 0.0187703
R9858 Y1.n786 Y1.n293 0.0187703
R9859 Y1.n789 Y1.n788 0.0187703
R9860 Y1.n814 Y1.n813 0.0187703
R9861 Y1.n821 Y1.n285 0.0187703
R9862 Y1.n824 Y1.n823 0.0187703
R9863 Y1.n829 Y1.n828 0.0187703
R9864 Y1.n832 Y1.n831 0.0187703
R9865 Y1.n841 Y1.n840 0.0187703
R9866 Y1.n845 Y1.n844 0.0187703
R9867 Y1.n849 Y1.n848 0.0187703
R9868 Y1.n851 Y1.n271 0.0187703
R9869 Y1.n860 Y1.n272 0.0187703
R9870 Y1.n276 Y1.n24 0.0187703
R9871 Y1.n1344 Y1.n26 0.0187703
R9872 Y1.n1202 Y1.n1201 0.0185541
R9873 Y1.n1323 Y1.n34 0.0185541
R9874 Y1.n464 Y1.n200 0.0185541
R9875 Y1.n673 Y1.n229 0.0185541
R9876 Y1.n976 Y1.n187 0.0184459
R9877 Y1.n1080 Y1.n1078 0.0184459
R9878 Y1.n734 Y1.n239 0.0184459
R9879 Y1.n810 Y1.n260 0.0184459
R9880 Y1.n1268 Y1.n1267 0.0182297
R9881 Y1.n572 Y1.n214 0.0182297
R9882 Y1.n977 Y1.n976 0.0181216
R9883 Y1.n1081 Y1.n1080 0.0181216
R9884 Y1.n734 Y1.n733 0.0181216
R9885 Y1.n810 Y1.n259 0.0181216
R9886 Y1.n71 Y1.n66 0.0175811
R9887 Y1.n1301 Y1.n10 0.0175811
R9888 Y1.n501 Y1.n500 0.0175811
R9889 Y1.n640 Y1.n223 0.0175811
R9890 Y1.n984 Y1.n983 0.0173649
R9891 Y1.n1095 Y1.n1094 0.0173649
R9892 Y1.n738 Y1.n240 0.0173649
R9893 Y1.n814 Y1.n261 0.0173649
R9894 Y1.n970 Y1.n969 0.0170405
R9895 Y1.n1084 Y1.n133 0.0170405
R9896 Y1.n307 Y1.n236 0.0170405
R9897 Y1.n806 Y1.n805 0.0170405
R9898 Y1.n1227 Y1.n61 0.0167162
R9899 Y1.n1287 Y1.n9 0.0167162
R9900 Y1.n523 Y1.n208 0.0167162
R9901 Y1.n618 Y1.n617 0.0167162
R9902 Y1.n994 Y1.n993 0.0162838
R9903 Y1.n1109 Y1.n119 0.0162838
R9904 Y1.n742 Y1.n241 0.0162838
R9905 Y1.n822 Y1.n821 0.0162838
R9906 Y1.n1372 Y1.n0 0.0161757
R9907 Y1.n1255 Y1.n1254 0.0159595
R9908 Y1.n1276 Y1.n4 0.0159595
R9909 Y1.n548 Y1.n213 0.0159595
R9910 Y1.n590 Y1.n361 0.0159595
R9911 Y1.n967 Y1.n189 0.0159595
R9912 Y1.n138 Y1.n132 0.0159595
R9913 Y1.n727 Y1.n235 0.0159595
R9914 Y1.n289 Y1.n256 0.0159595
R9915 Y1.n1190 Y1.n1189 0.0157432
R9916 Y1.n1332 Y1.n18 0.0157432
R9917 Y1.n440 Y1.n199 0.0157432
R9918 Y1.n698 Y1.n230 0.0157432
R9919 Y1.n80 Y1.n75 0.0152027
R9920 Y1.n1319 Y1.n15 0.0152027
R9921 Y1.n473 Y1.n404 0.0152027
R9922 Y1.n665 Y1.n228 0.0152027
R9923 Y1.n1002 Y1.n173 0.0152027
R9924 Y1.n1101 Y1.n120 0.0152027
R9925 Y1.n748 Y1.n747 0.0152027
R9926 Y1.n824 Y1.n264 0.0152027
R9927 Y1.n1272 Y1.n3 0.0148784
R9928 Y1.n581 Y1.n215 0.0148784
R9929 Y1.n958 Y1.n957 0.0148784
R9930 Y1.n1068 Y1.n1067 0.0148784
R9931 Y1.n723 Y1.n234 0.0148784
R9932 Y1.n796 Y1.n255 0.0148784
R9933 Y1.n1221 Y1.n70 0.0141216
R9934 Y1.n1305 Y1.n1303 0.0141216
R9935 Y1.n489 Y1.n205 0.0141216
R9936 Y1.n647 Y1.n224 0.0141216
R9937 Y1.n174 Y1.n167 0.0141216
R9938 Y1.n1119 Y1.n115 0.0141216
R9939 Y1.n750 Y1.n244 0.0141216
R9940 Y1.n829 Y1.n265 0.0141216
R9941 Y1.n1180 Y1.n1179 0.0137973
R9942 Y1.n1178 Y1.n90 0.0137973
R9943 Y1.n1056 Y1.n1055 0.0137973
R9944 Y1.n1177 Y1.n89 0.0137973
R9945 Y1.n792 Y1.n254 0.0137973
R9946 Y1.n25 Y1.n21 0.0137973
R9947 Y1.n1350 Y1.n20 0.0137973
R9948 Y1.n1349 Y1.n1348 0.0137973
R9949 Y1.n855 Y1.n30 0.0134381
R9950 Y1.n1241 Y1.n1240 0.0133649
R9951 Y1.n1285 Y1.n8 0.0133649
R9952 Y1.n530 Y1.n209 0.0133649
R9953 Y1.n606 Y1.n220 0.0133649
R9954 Y1.n1019 Y1.n1018 0.0130405
R9955 Y1.n1120 Y1.n111 0.0130405
R9956 Y1.n752 Y1.n245 0.0130405
R9957 Y1.n831 Y1.n266 0.0130405
R9958 Y1.n1058 Y1.n1054 0.0128243
R9959 Y1.n1166 Y1.n93 0.0128243
R9960 Y1.n788 Y1.n787 0.0128243
R9961 Y1.n1345 Y1.n1344 0.0128243
R9962 Y1.n59 Y1.n58 0.0126081
R9963 Y1.n44 Y1.n5 0.0126081
R9964 Y1.n547 Y1.n546 0.0126081
R9965 Y1.n599 Y1.n218 0.0126081
R9966 Y1.n1184 Y1.n1183 0.0123919
R9967 Y1.n28 Y1.n19 0.0123919
R9968 Y1.n434 Y1.n198 0.0123919
R9969 Y1.n712 Y1.n320 0.0123919
R9970 Y1.n1015 Y1.n1011 0.0119595
R9971 Y1.n1129 Y1.n108 0.0119595
R9972 Y1.n763 Y1.n246 0.0119595
R9973 Y1.n841 Y1.n281 0.0119595
R9974 Y1.n1208 Y1.n73 0.0118514
R9975 Y1.n1315 Y1.n14 0.0118514
R9976 Y1.n482 Y1.n203 0.0118514
R9977 Y1.n664 Y1.n663 0.0118514
R9978 Y1.n1038 Y1.n1037 0.0117432
R9979 Y1.n1165 Y1.n1164 0.0117432
R9980 Y1.n293 Y1.n251 0.0117432
R9981 Y1.n276 Y1.n275 0.0117432
R9982 Y1.n1172 Y1.n1171 0.0116588
R9983 Y1.n1184 Y1.n89 0.011527
R9984 Y1.n434 Y1.n433 0.011527
R9985 Y1.n28 Y1.n21 0.0114189
R9986 Y1.n715 Y1.n712 0.0114189
R9987 Y1.n313 Y1.n312 0.0109762
R9988 Y1.n311 Y1.n310 0.0109762
R9989 Y1.n756 Y1.n301 0.0109762
R9990 Y1.n759 Y1.n758 0.0109762
R9991 Y1.n757 Y1.n295 0.0109762
R9992 Y1.n783 Y1.n782 0.0109762
R9993 Y1.n800 Y1.n291 0.0109762
R9994 Y1.n801 Y1.n287 0.0109762
R9995 Y1.n818 Y1.n817 0.0109762
R9996 Y1.n835 Y1.n283 0.0109762
R9997 Y1.n837 Y1.n836 0.0109762
R9998 Y1.n854 Y1.n278 0.0109762
R9999 Y1.n856 Y1.n855 0.0109762
R10000 Y1.n1195 Y1.n85 0.0109762
R10001 Y1.n1198 Y1.n1195 0.0109762
R10002 Y1.n1198 Y1.n1197 0.0109762
R10003 Y1.n1197 Y1.n1196 0.0109762
R10004 Y1.n1196 Y1.n63 0.0109762
R10005 Y1.n1233 Y1.n63 0.0109762
R10006 Y1.n1235 Y1.n1233 0.0109762
R10007 Y1.n1235 Y1.n1234 0.0109762
R10008 Y1.n1234 Y1.n50 0.0109762
R10009 Y1.n1258 Y1.n50 0.0109762
R10010 Y1.n1262 Y1.n1258 0.0109762
R10011 Y1.n1261 Y1.n1260 0.0109762
R10012 Y1.n1260 Y1.n1259 0.0109762
R10013 Y1.n1259 Y1.n42 0.0109762
R10014 Y1.n1291 Y1.n42 0.0109762
R10015 Y1.n1292 Y1.n1291 0.0109762
R10016 Y1.n1292 Y1.n38 0.0109762
R10017 Y1.n1308 Y1.n38 0.0109762
R10018 Y1.n1311 Y1.n1308 0.0109762
R10019 Y1.n1311 Y1.n1310 0.0109762
R10020 Y1.n1310 Y1.n1309 0.0109762
R10021 Y1.n1309 Y1.n32 0.0109762
R10022 Y1.n1336 Y1.n32 0.0109762
R10023 Y1.n964 Y1.n180 0.0109762
R10024 Y1.n990 Y1.n989 0.0109762
R10025 Y1.n1023 Y1.n164 0.0109762
R10026 Y1.n1025 Y1.n1024 0.0109762
R10027 Y1.n1026 Y1.n156 0.0109762
R10028 Y1.n1061 Y1.n147 0.0109762
R10029 Y1.n1062 Y1.n129 0.0109762
R10030 Y1.n1089 Y1.n1088 0.0109762
R10031 Y1.n1090 Y1.n121 0.0109762
R10032 Y1.n1124 Y1.n113 0.0109762
R10033 Y1.n1125 Y1.n106 0.0109762
R10034 Y1.n312 Y1.n311 0.01095
R10035 Y1.n310 Y1.n301 0.01095
R10036 Y1.n759 Y1.n756 0.01095
R10037 Y1.n758 Y1.n757 0.01095
R10038 Y1.n782 Y1.n295 0.01095
R10039 Y1.n783 Y1.n291 0.01095
R10040 Y1.n801 Y1.n800 0.01095
R10041 Y1.n817 Y1.n287 0.01095
R10042 Y1.n818 Y1.n283 0.01095
R10043 Y1.n837 Y1.n835 0.01095
R10044 Y1.n836 Y1.n278 0.01095
R10045 Y1.n856 Y1.n854 0.01095
R10046 Y1.n1262 Y1.n1261 0.01095
R10047 Y1.n1337 Y1.n1336 0.01095
R10048 Y1.n964 Y1.n963 0.01095
R10049 Y1.n989 Y1.n180 0.01095
R10050 Y1.n990 Y1.n164 0.01095
R10051 Y1.n1024 Y1.n1023 0.01095
R10052 Y1.n1026 Y1.n1025 0.01095
R10053 Y1.n156 Y1.n147 0.01095
R10054 Y1.n1062 Y1.n1061 0.01095
R10055 Y1.n1088 Y1.n129 0.01095
R10056 Y1.n1090 Y1.n1089 0.01095
R10057 Y1.n121 Y1.n113 0.01095
R10058 Y1.n1125 Y1.n1124 0.01095
R10059 Y1.n1139 Y1.n106 0.01095
R10060 Y1.n1012 Y1.n158 0.0108784
R10061 Y1.n1135 Y1.n1134 0.0108784
R10062 Y1.n767 Y1.n298 0.0108784
R10063 Y1.n845 Y1.n269 0.0108784
R10064 Y1.n1214 Y1.n1213 0.0107703
R10065 Y1.n1314 Y1.n13 0.0107703
R10066 Y1.n483 Y1.n204 0.0107703
R10067 Y1.n336 Y1.n225 0.0107703
R10068 Y1.n1048 Y1.n1047 0.0106622
R10069 Y1.n1143 Y1.n1142 0.0106622
R10070 Y1.n778 Y1.n250 0.0106622
R10071 Y1.n861 Y1.n860 0.0106622
R10072 Y1.n1171 Y1.n85 0.0106095
R10073 Y1.n1248 Y1.n1247 0.0100135
R10074 Y1.n1283 Y1.n1282 0.0100135
R10075 Y1.n379 Y1.n210 0.0100135
R10076 Y1.n600 Y1.n219 0.0100135
R10077 Y1.n1031 Y1.n1030 0.0097973
R10078 Y1.n1158 Y1.n102 0.0097973
R10079 Y1.n771 Y1.n249 0.0097973
R10080 Y1.n849 Y1.n270 0.0097973
R10081 Y1.n1173 Y1.n1172 0.00967266
R10082 Y1.n1032 Y1.n1031 0.00958108
R10083 Y1.n1158 Y1.n1157 0.00958108
R10084 Y1.n774 Y1.n249 0.00958108
R10085 Y1.n851 Y1.n270 0.00958108
R10086 Y1.n1248 Y1.n57 0.00925676
R10087 Y1.n1284 Y1.n1283 0.00925676
R10088 Y1.n531 Y1.n210 0.00925676
R10089 Y1.n607 Y1.n219 0.00925676
R10090 Y1.n1041 Y1.n147 0.00880612
R10091 Y1.n1048 Y1.n154 0.00871622
R10092 Y1.n1142 Y1.n103 0.00871622
R10093 Y1.n775 Y1.n250 0.00871622
R10094 Y1.n861 Y1.n271 0.00871622
R10095 Y1.n1215 Y1.n1214 0.0085
R10096 Y1.n1304 Y1.n13 0.0085
R10097 Y1.n490 Y1.n204 0.0085
R10098 Y1.n648 Y1.n225 0.0085
R10099 Y1.n1029 Y1.n158 0.0085
R10100 Y1.n1136 Y1.n1135 0.0085
R10101 Y1.n770 Y1.n298 0.0085
R10102 Y1.n848 Y1.n269 0.0085
R10103 Y1.n314 Y1.n313 0.00809524
R10104 Y1.n1170 Y1.n96 0.00778095
R10105 Y1.n1037 Y1.n155 0.00763514
R10106 Y1.n1164 Y1.n98 0.00763514
R10107 Y1.n779 Y1.n251 0.00763514
R10108 Y1.n275 Y1.n272 0.00763514
R10109 Y1.n1209 Y1.n1208 0.00741892
R10110 Y1.n1318 Y1.n14 0.00741892
R10111 Y1.n474 Y1.n203 0.00741892
R10112 Y1.n666 Y1.n664 0.00741892
R10113 Y1.n1015 Y1.n1014 0.00741892
R10114 Y1.n1133 Y1.n108 0.00741892
R10115 Y1.n766 Y1.n246 0.00741892
R10116 Y1.n844 Y1.n281 0.00741892
R10117 Y1.n1154 Y1.n1139 0.00725714
R10118 Y1.n1173 Y1.n1170 0.00707381
R10119 Y1.n1183 Y1.n87 0.00698649
R10120 Y1.n1333 Y1.n19 0.00698649
R10121 Y1.n441 Y1.n198 0.00698649
R10122 Y1.n699 Y1.n320 0.00698649
R10123 Y1.n963 Y1.n193 0.00696162
R10124 Y1.n1339 Y1.n1337 0.00691667
R10125 Y1.n58 Y1.n52 0.00666216
R10126 Y1.n1277 Y1.n5 0.00666216
R10127 Y1.n549 Y1.n547 0.00666216
R10128 Y1.n591 Y1.n218 0.00666216
R10129 Y1.n1054 Y1.n150 0.00655405
R10130 Y1.n1167 Y1.n1166 0.00655405
R10131 Y1.n787 Y1.n786 0.00655405
R10132 Y1.n1345 Y1.n24 0.00655405
R10133 Y1.n1018 Y1.n169 0.00633784
R10134 Y1.n1128 Y1.n111 0.00633784
R10135 Y1.n762 Y1.n245 0.00633784
R10136 Y1.n840 Y1.n266 0.00633784
R10137 Y1.n1240 Y1.n1239 0.00590541
R10138 Y1.n1288 Y1.n8 0.00590541
R10139 Y1.n524 Y1.n209 0.00590541
R10140 Y1.n616 Y1.n220 0.00590541
R10141 Y1.n142 Y1.n129 0.00588776
R10142 Y1.n963 Y1.n192 0.00588776
R10143 Y1.n1057 Y1.n1056 0.00547297
R10144 Y1.n1177 Y1.n1176 0.00547297
R10145 Y1.n789 Y1.n254 0.00547297
R10146 Y1.n26 Y1.n25 0.00547297
R10147 Y1.n1020 Y1.n167 0.00525676
R10148 Y1.n1121 Y1.n1119 0.00525676
R10149 Y1.n753 Y1.n244 0.00525676
R10150 Y1.n832 Y1.n265 0.00525676
R10151 Y1.n1221 Y1.n1220 0.00514865
R10152 Y1.n1303 Y1.n1302 0.00514865
R10153 Y1.n499 Y1.n205 0.00514865
R10154 Y1.n641 Y1.n224 0.00514865
R10155 Y1.n1338 Y1.n30 0.00440238
R10156 Y1.n1269 Y1.n3 0.00439189
R10157 Y1.n573 Y1.n215 0.00439189
R10158 Y1.n957 Y1.n195 0.00439189
R10159 Y1.n1068 Y1.n137 0.00439189
R10160 Y1.n714 Y1.n234 0.00439189
R10161 Y1.n793 Y1.n255 0.00439189
R10162 Y1.n1186 Y1.n1185 0.00425921
R10163 Y1.n1188 Y1.n86 0.00425921
R10164 Y1.n1212 Y1.n1211 0.00425921
R10165 Y1.n1217 Y1.n1216 0.00425921
R10166 Y1.n65 Y1.n62 0.00425921
R10167 Y1.n1238 Y1.n1237 0.00425921
R10168 Y1.n1243 Y1.n1242 0.00425921
R10169 Y1.n1246 Y1.n1245 0.00425921
R10170 Y1.n1270 Y1.n47 0.00425921
R10171 Y1.n1281 Y1.n1279 0.00425921
R10172 Y1.n1286 Y1.n43 0.00425921
R10173 Y1.n1289 Y1.n41 0.00425921
R10174 Y1.n1294 Y1.n40 0.00425921
R10175 Y1.n1306 Y1.n37 0.00425921
R10176 Y1.n1316 Y1.n1313 0.00425921
R10177 Y1.n1331 Y1.n1330 0.00425921
R10178 Y1.n1334 Y1.n29 0.00425921
R10179 Y1.n1028 Y1.n159 0.00425921
R10180 Y1.n1033 Y1.n157 0.00425921
R10181 Y1.n1137 Y1.n107 0.00425921
R10182 Y1.n1156 Y1.n104 0.00425921
R10183 Y1.n731 Y1.n730 0.00425921
R10184 Y1.n736 Y1.n735 0.00425921
R10185 Y1.n740 Y1.n739 0.00425921
R10186 Y1.n744 Y1.n743 0.00425921
R10187 Y1.n765 Y1.n764 0.00425921
R10188 Y1.n769 Y1.n768 0.00425921
R10189 Y1.n773 Y1.n772 0.00425921
R10190 Y1.n777 Y1.n776 0.00425921
R10191 Y1.n794 Y1.n791 0.00425921
R10192 Y1.n808 Y1.n288 0.00425921
R10193 Y1.n812 Y1.n811 0.00425921
R10194 Y1.n815 Y1.n286 0.00425921
R10195 Y1.n820 Y1.n284 0.00425921
R10196 Y1.n843 Y1.n842 0.00425921
R10197 Y1.n847 Y1.n846 0.00425921
R10198 Y1.n852 Y1.n850 0.00425921
R10199 Y1.n859 Y1.n273 0.00425921
R10200 Y1.n1152 Y1.n1151 0.00424524
R10201 Y1.n1193 Y1.n86 0.0042371
R10202 Y1.n1200 Y1.n82 0.0042371
R10203 Y1.n84 Y1.n83 0.0042371
R10204 Y1.n1211 Y1.n1210 0.0042371
R10205 Y1.n1219 Y1.n64 0.0042371
R10206 Y1.n1231 Y1.n65 0.0042371
R10207 Y1.n1245 Y1.n51 0.0042371
R10208 Y1.n1256 Y1.n49 0.0042371
R10209 Y1.n1265 Y1.n1264 0.0042371
R10210 Y1.n1265 Y1.n47 0.0042371
R10211 Y1.n1271 Y1.n1270 0.0042371
R10212 Y1.n1275 Y1.n1274 0.0042371
R10213 Y1.n1279 Y1.n1278 0.0042371
R10214 Y1.n1298 Y1.n40 0.0042371
R10215 Y1.n1300 Y1.n39 0.0042371
R10216 Y1.n1317 Y1.n1316 0.0042371
R10217 Y1.n1321 Y1.n1320 0.0042371
R10218 Y1.n1326 Y1.n1324 0.0042371
R10219 Y1.n1330 Y1.n33 0.0042371
R10220 Y1.n971 Y1.n188 0.0042371
R10221 Y1.n1000 Y1.n165 0.0042371
R10222 Y1.n1021 Y1.n166 0.0042371
R10223 Y1.n1059 Y1.n149 0.0042371
R10224 Y1.n1086 Y1.n131 0.0042371
R10225 Y1.n1103 Y1.n114 0.0042371
R10226 Y1.n1122 Y1.n112 0.0042371
R10227 Y1.n1168 Y1.n97 0.0042371
R10228 Y1.n1175 Y1.n94 0.0042371
R10229 Y1.n726 Y1.n725 0.0042371
R10230 Y1.n730 Y1.n729 0.0042371
R10231 Y1.n746 Y1.n744 0.0042371
R10232 Y1.n751 Y1.n302 0.0042371
R10233 Y1.n754 Y1.n300 0.0042371
R10234 Y1.n764 Y1.n761 0.0042371
R10235 Y1.n780 Y1.n777 0.0042371
R10236 Y1.n785 Y1.n294 0.0042371
R10237 Y1.n790 Y1.n292 0.0042371
R10238 Y1.n791 Y1.n790 0.0042371
R10239 Y1.n795 Y1.n794 0.0042371
R10240 Y1.n798 Y1.n290 0.0042371
R10241 Y1.n803 Y1.n288 0.0042371
R10242 Y1.n825 Y1.n284 0.0042371
R10243 Y1.n830 Y1.n827 0.0042371
R10244 Y1.n833 Y1.n282 0.0042371
R10245 Y1.n842 Y1.n839 0.0042371
R10246 Y1.n859 Y1.n858 0.0042371
R10247 Y1.n277 Y1.n274 0.0042371
R10248 Y1.n1343 Y1.n1342 0.0042371
R10249 Y1.n1342 Y1.n1341 0.0042371
R10250 Y1.n718 Y1.n717 0.00423273
R10251 Y1.n429 Y1.n428 0.00422178
R10252 Y1.n705 Y1.n317 0.00422178
R10253 Y1.n1154 Y1.n1153 0.00421905
R10254 Y1.n1002 Y1.n1001 0.00417568
R10255 Y1.n1102 Y1.n1101 0.00417568
R10256 Y1.n749 Y1.n748 0.00417568
R10257 Y1.n828 Y1.n264 0.00417568
R10258 Y1.n1194 Y1.n82 0.00410442
R10259 Y1.n1326 Y1.n1325 0.00410442
R10260 Y1.n81 Y1.n80 0.00406757
R10261 Y1.n1322 Y1.n15 0.00406757
R10262 Y1.n465 Y1.n404 0.00406757
R10263 Y1.n674 Y1.n228 0.00406757
R10264 Y1.n1040 Y1.n148 0.00402269
R10265 Y1.n975 Y1.n178 0.00398793
R10266 Y1.n1079 Y1.n126 0.00398793
R10267 Y1.n735 Y1.n306 0.00397174
R10268 Y1.n773 Y1.n296 0.00397174
R10269 Y1.n811 Y1.n809 0.00397174
R10270 Y1.n853 Y1.n852 0.00397174
R10271 Y1.n1244 Y1.n1243 0.00394963
R10272 Y1.n1280 Y1.n43 0.00394963
R10273 Y1.n966 Y1.n190 0.00394626
R10274 Y1.n141 Y1.n130 0.00394626
R10275 Y1.n421 Y1.n191 0.00393696
R10276 Y1.n1065 Y1.n1064 0.00393696
R10277 Y1.n985 Y1.n177 0.00390294
R10278 Y1.n1097 Y1.n122 0.00390294
R10279 Y1.n1046 Y1.n1045 0.00389381
R10280 Y1.n996 Y1.n175 0.00385851
R10281 Y1.n1010 Y1.n160 0.00385851
R10282 Y1.n1107 Y1.n1100 0.00385851
R10283 Y1.n1131 Y1.n1130 0.00385851
R10284 Y1.n997 Y1.n996 0.00380768
R10285 Y1.n1107 Y1.n1106 0.00380768
R10286 Y1.n1010 Y1.n163 0.00380053
R10287 Y1.n1130 Y1.n110 0.00380053
R10288 Y1.n1216 Y1.n72 0.00379484
R10289 Y1.n1312 Y1.n37 0.00379484
R10290 Y1.n716 Y1.n316 0.00379484
R10291 Y1.n1174 Y1.n95 0.00377273
R10292 Y1.n972 Y1.n971 0.0037725
R10293 Y1.n1046 Y1.n1036 0.0037725
R10294 Y1.n131 Y1.n127 0.0037725
R10295 Y1.n1150 Y1.n1149 0.00374762
R10296 Y1.n1064 Y1.n1063 0.00372958
R10297 Y1.n745 Y1.n302 0.0037285
R10298 Y1.n827 Y1.n826 0.0037285
R10299 Y1.n149 Y1.n146 0.00372177
R10300 Y1.n760 Y1.n300 0.00370639
R10301 Y1.n838 Y1.n282 0.00370639
R10302 Y1.n1148 Y1.n96 0.00369524
R10303 Y1.n1232 Y1.n64 0.00366216
R10304 Y1.n1300 Y1.n1299 0.00366216
R10305 Y1.n1141 Y1.n1140 0.00366216
R10306 Y1.n1155 Y1.n105 0.00364005
R10307 Y1.n1191 Y1.n1190 0.00363514
R10308 Y1.n1329 Y1.n18 0.00363514
R10309 Y1.n411 Y1.n199 0.00363514
R10310 Y1.n690 Y1.n230 0.00363514
R10311 Y1.n721 Y1.n719 0.00359048
R10312 Y1.n1034 Y1.n1033 0.00358532
R10313 Y1.n428 Y1.n424 0.00357902
R10314 Y1.n705 Y1.n704 0.00357902
R10315 Y1.n975 Y1.n974 0.00357098
R10316 Y1.n1079 Y1.n128 0.00357098
R10317 Y1.n1237 Y1.n1236 0.00348526
R10318 Y1.n1293 Y1.n41 0.00348526
R10319 Y1.n1000 Y1.n999 0.003457
R10320 Y1.n1104 Y1.n1103 0.003457
R10321 Y1.n166 Y1.n162 0.00344926
R10322 Y1.n1126 Y1.n112 0.00344926
R10323 Y1.n740 Y1.n304 0.00344103
R10324 Y1.n768 Y1.n299 0.00344103
R10325 Y1.n819 Y1.n286 0.00344103
R10326 Y1.n846 Y1.n280 0.00344103
R10327 Y1.n1013 Y1.n161 0.00343273
R10328 Y1.n1132 Y1.n109 0.00343273
R10329 Y1.n992 Y1.n991 0.00341839
R10330 Y1.n1099 Y1.n1098 0.00341839
R10331 Y1.n1091 Y1.n1090 0.00341837
R10332 Y1.n989 Y1.n179 0.00341837
R10333 Y1.n720 Y1.n314 0.00335476
R10334 Y1.n83 Y1.n74 0.00335258
R10335 Y1.n1320 Y1.n36 0.00335258
R10336 Y1.n991 Y1.n177 0.0033136
R10337 Y1.n1098 Y1.n1097 0.0033136
R10338 Y1.n1254 Y1.n53 0.00331081
R10339 Y1.n1273 Y1.n4 0.00331081
R10340 Y1.n372 Y1.n213 0.00331081
R10341 Y1.n582 Y1.n361 0.00331081
R10342 Y1.n959 Y1.n189 0.00331081
R10343 Y1.n139 Y1.n138 0.00331081
R10344 Y1.n724 Y1.n235 0.00331081
R10345 Y1.n797 Y1.n256 0.00331081
R10346 Y1.n168 Y1.n162 0.00330444
R10347 Y1.n1127 Y1.n1126 0.00330444
R10348 Y1.n161 Y1.n159 0.0032992
R10349 Y1.n109 Y1.n107 0.0032992
R10350 Y1.n999 Y1.n998 0.00329663
R10351 Y1.n1105 Y1.n1104 0.00329663
R10352 Y1.n1146 Y1.n1145 0.00324201
R10353 Y1.n1257 Y1.n1256 0.00319779
R10354 Y1.n1275 Y1.n45 0.00319779
R10355 Y1.n1147 Y1.n97 0.00319779
R10356 Y1.n781 Y1.n294 0.00319779
R10357 Y1.n857 Y1.n277 0.00319779
R10358 Y1.n966 Y1.n965 0.00317568
R10359 Y1.n1087 Y1.n130 0.00317568
R10360 Y1.n726 Y1.n308 0.00317568
R10361 Y1.n802 Y1.n290 0.00317568
R10362 Y1.n974 Y1.n973 0.00316007
R10363 Y1.n1076 Y1.n128 0.00316007
R10364 Y1.n1035 Y1.n1034 0.00314581
R10365 Y1.n722 Y1.n315 0.00310934
R10366 Y1.n995 Y1.n994 0.00309459
R10367 Y1.n1109 Y1.n1108 0.00309459
R10368 Y1.n303 Y1.n241 0.00309459
R10369 Y1.n823 Y1.n822 0.00309459
R10370 Y1.n1187 Y1.n1186 0.003043
R10371 Y1.n1335 Y1.n1334 0.003043
R10372 Y1.n1063 Y1.n145 0.00302306
R10373 Y1.n146 Y1.n145 0.00300884
R10374 Y1.n470 Y1.n468 0.0029881
R10375 Y1.n505 Y1.n504 0.0029881
R10376 Y1.n520 Y1.n386 0.0029881
R10377 Y1.n622 Y1.n621 0.0029881
R10378 Y1.n1036 Y1.n1035 0.00298054
R10379 Y1.n973 Y1.n972 0.00298054
R10380 Y1.n1076 Y1.n127 0.00298054
R10381 Y1.n637 Y1.n343 0.0029619
R10382 Y1.n671 Y1.n670 0.0029619
R10383 Y1.n168 Y1.n163 0.00293083
R10384 Y1.n1127 Y1.n110 0.00293083
R10385 Y1.n998 Y1.n997 0.0029237
R10386 Y1.n1106 Y1.n1105 0.0029237
R10387 Y1.n1263 Y1.n49 0.00291032
R10388 Y1.n1274 Y1.n46 0.00291032
R10389 Y1.n1060 Y1.n148 0.00291032
R10390 Y1.n1169 Y1.n1168 0.00291032
R10391 Y1.n725 Y1.n309 0.00291032
R10392 Y1.n785 Y1.n784 0.00291032
R10393 Y1.n799 Y1.n798 0.00291032
R10394 Y1.n274 Y1.n27 0.00291032
R10395 Y1.n992 Y1.n175 0.00289527
R10396 Y1.n1100 Y1.n1099 0.00289527
R10397 Y1.n1013 Y1.n160 0.00289527
R10398 Y1.n1132 Y1.n1131 0.00289527
R10399 Y1.n426 Y1.n424 0.00287188
R10400 Y1.n707 Y1.n704 0.00284569
R10401 Y1.n1045 Y1.n1044 0.00283826
R10402 Y1.n1339 Y1.n1338 0.00283095
R10403 Y1.n194 Y1.n191 0.00279542
R10404 Y1.n1066 Y1.n1065 0.00279542
R10405 Y1.n181 Y1.n178 0.00276679
R10406 Y1.n126 Y1.n125 0.00276679
R10407 Y1.n1199 Y1.n84 0.00275553
R10408 Y1.n1321 Y1.n35 0.00275553
R10409 Y1.n1185 Y1.n88 0.00273342
R10410 Y1.n1341 Y1.n29 0.00273342
R10411 Y1.n426 Y1.n425 0.00272619
R10412 Y1.n425 Y1.n418 0.00272619
R10413 Y1.n444 Y1.n416 0.00272619
R10414 Y1.n446 Y1.n445 0.00272619
R10415 Y1.n454 Y1.n453 0.00272619
R10416 Y1.n462 Y1.n406 0.00272619
R10417 Y1.n467 Y1.n406 0.00272619
R10418 Y1.n469 Y1.n402 0.00272619
R10419 Y1.n477 Y1.n402 0.00272619
R10420 Y1.n485 Y1.n399 0.00272619
R10421 Y1.n486 Y1.n485 0.00272619
R10422 Y1.n495 Y1.n494 0.00272619
R10423 Y1.n496 Y1.n495 0.00272619
R10424 Y1.n506 Y1.n393 0.00272619
R10425 Y1.n510 Y1.n393 0.00272619
R10426 Y1.n518 Y1.n389 0.00272619
R10427 Y1.n519 Y1.n518 0.00272619
R10428 Y1.n527 Y1.n526 0.00272619
R10429 Y1.n528 Y1.n383 0.00272619
R10430 Y1.n540 Y1.n381 0.00272619
R10431 Y1.n552 Y1.n377 0.00272619
R10432 Y1.n553 Y1.n552 0.00272619
R10433 Y1.n559 Y1.n558 0.00272619
R10434 Y1.n561 Y1.n559 0.00272619
R10435 Y1.n561 Y1.n560 0.00272619
R10436 Y1.n570 Y1.n569 0.00272619
R10437 Y1.n579 Y1.n578 0.00272619
R10438 Y1.n578 Y1.n363 0.00272619
R10439 Y1.n588 Y1.n587 0.00272619
R10440 Y1.n587 Y1.n359 0.00272619
R10441 Y1.n594 Y1.n359 0.00272619
R10442 Y1.n602 Y1.n356 0.00272619
R10443 Y1.n603 Y1.n602 0.00272619
R10444 Y1.n612 Y1.n611 0.00272619
R10445 Y1.n613 Y1.n612 0.00272619
R10446 Y1.n627 Y1.n350 0.00272619
R10447 Y1.n636 Y1.n635 0.00272619
R10448 Y1.n644 Y1.n643 0.00272619
R10449 Y1.n645 Y1.n340 0.00272619
R10450 Y1.n657 Y1.n338 0.00272619
R10451 Y1.n669 Y1.n334 0.00272619
R10452 Y1.n670 Y1.n669 0.00272619
R10453 Y1.n677 Y1.n332 0.00272619
R10454 Y1.n678 Y1.n677 0.00272619
R10455 Y1.n679 Y1.n678 0.00272619
R10456 Y1.n687 Y1.n685 0.00272619
R10457 Y1.n687 Y1.n686 0.00272619
R10458 Y1.n696 Y1.n694 0.00272619
R10459 Y1.n696 Y1.n695 0.00272619
R10460 Y1.n710 Y1.n709 0.00272619
R10461 Y1.n708 Y1.n707 0.00272619
R10462 Y1.n436 Y1.n418 0.0027
R10463 Y1.n445 Y1.n444 0.0027
R10464 Y1.n454 Y1.n452 0.0027
R10465 Y1.n462 Y1.n461 0.0027
R10466 Y1.n470 Y1.n469 0.0027
R10467 Y1.n496 Y1.n395 0.0027
R10468 Y1.n528 Y1.n527 0.0027
R10469 Y1.n536 Y1.n381 0.0027
R10470 Y1.n542 Y1.n377 0.0027
R10471 Y1.n570 Y1.n568 0.0027
R10472 Y1.n579 Y1.n577 0.0027
R10473 Y1.n613 Y1.n352 0.0027
R10474 Y1.n623 Y1.n350 0.0027
R10475 Y1.n635 Y1.n346 0.0027
R10476 Y1.n645 Y1.n644 0.0027
R10477 Y1.n653 Y1.n338 0.0027
R10478 Y1.n659 Y1.n334 0.0027
R10479 Y1.n695 Y1.n322 0.0027
R10480 Y1.n709 Y1.n708 0.0027
R10481 Y1.n504 Y1.n395 0.00264762
R10482 Y1.n643 Y1.n343 0.00264762
R10483 Y1.n739 Y1.n305 0.00264496
R10484 Y1.n816 Y1.n815 0.00264496
R10485 Y1.n1028 Y1.n1027 0.00262285
R10486 Y1.n1138 Y1.n1137 0.00262285
R10487 Y1.n769 Y1.n297 0.00262285
R10488 Y1.n847 Y1.n279 0.00262285
R10489 Y1.n520 Y1.n519 0.00262143
R10490 Y1.n623 Y1.n622 0.00262143
R10491 Y1.n1238 Y1.n60 0.00260074
R10492 Y1.n1290 Y1.n1289 0.00260074
R10493 Y1.n472 Y1.n405 0.00257862
R10494 Y1.n672 Y1.n333 0.00257862
R10495 Y1.n621 Y1.n352 0.00256905
R10496 Y1.n1228 Y1.n1227 0.00255405
R10497 Y1.n1295 Y1.n9 0.00255405
R10498 Y1.n516 Y1.n208 0.00255405
R10499 Y1.n617 Y1.n348 0.00255405
R10500 Y1.n526 Y1.n386 0.00254286
R10501 Y1.n637 Y1.n636 0.00254286
R10502 Y1.n522 Y1.n387 0.0025344
R10503 Y1.n506 Y1.n505 0.00251667
R10504 Y1.n620 Y1.n619 0.00251228
R10505 Y1.n431 Y1.n430 0.0024936
R10506 Y1.n468 Y1.n467 0.00246429
R10507 Y1.n671 Y1.n332 0.00246429
R10508 Y1.n1219 Y1.n1218 0.00244595
R10509 Y1.n1307 Y1.n39 0.00244595
R10510 Y1.n487 Y1.n486 0.0024381
R10511 Y1.n653 Y1.n652 0.0024381
R10512 Y1.n503 Y1.n502 0.00242383
R10513 Y1.n639 Y1.n344 0.00242383
R10514 Y1.n719 Y1.n718 0.00238571
R10515 Y1.n1151 Y1.n1150 0.00238571
R10516 Y1.n451 Y1.n414 0.00238571
R10517 Y1.n460 Y1.n409 0.00238571
R10518 Y1.n479 Y1.n478 0.00238571
R10519 Y1.n487 Y1.n397 0.00238571
R10520 Y1.n512 Y1.n511 0.00238571
R10521 Y1.n535 Y1.n534 0.00238571
R10522 Y1.n543 Y1.n541 0.00238571
R10523 Y1.n567 Y1.n370 0.00238571
R10524 Y1.n576 Y1.n366 0.00238571
R10525 Y1.n585 Y1.n363 0.00238571
R10526 Y1.n596 Y1.n595 0.00238571
R10527 Y1.n604 Y1.n354 0.00238571
R10528 Y1.n629 Y1.n628 0.00238571
R10529 Y1.n652 Y1.n651 0.00238571
R10530 Y1.n660 Y1.n658 0.00238571
R10531 Y1.n684 Y1.n330 0.00238571
R10532 Y1.n693 Y1.n325 0.00238571
R10533 Y1.n443 Y1.n442 0.00237961
R10534 Y1.n447 Y1.n415 0.00237961
R10535 Y1.n455 Y1.n413 0.00237961
R10536 Y1.n463 Y1.n407 0.00237961
R10537 Y1.n466 Y1.n407 0.00237961
R10538 Y1.n475 Y1.n403 0.00237961
R10539 Y1.n476 Y1.n475 0.00237961
R10540 Y1.n484 Y1.n400 0.00237961
R10541 Y1.n484 Y1.n398 0.00237961
R10542 Y1.n493 Y1.n396 0.00237961
R10543 Y1.n497 Y1.n396 0.00237961
R10544 Y1.n508 Y1.n507 0.00237961
R10545 Y1.n509 Y1.n508 0.00237961
R10546 Y1.n517 Y1.n390 0.00237961
R10547 Y1.n517 Y1.n388 0.00237961
R10548 Y1.n525 Y1.n385 0.00237961
R10549 Y1.n529 Y1.n384 0.00237961
R10550 Y1.n539 Y1.n538 0.00237961
R10551 Y1.n551 Y1.n550 0.00237961
R10552 Y1.n551 Y1.n376 0.00237961
R10553 Y1.n557 Y1.n373 0.00237961
R10554 Y1.n562 Y1.n373 0.00237961
R10555 Y1.n562 Y1.n374 0.00237961
R10556 Y1.n571 Y1.n369 0.00237961
R10557 Y1.n580 Y1.n364 0.00237961
R10558 Y1.n583 Y1.n364 0.00237961
R10559 Y1.n589 Y1.n360 0.00237961
R10560 Y1.n592 Y1.n360 0.00237961
R10561 Y1.n593 Y1.n592 0.00237961
R10562 Y1.n601 Y1.n357 0.00237961
R10563 Y1.n601 Y1.n355 0.00237961
R10564 Y1.n610 Y1.n353 0.00237961
R10565 Y1.n614 Y1.n353 0.00237961
R10566 Y1.n626 Y1.n625 0.00237961
R10567 Y1.n634 Y1.n345 0.00237961
R10568 Y1.n642 Y1.n342 0.00237961
R10569 Y1.n646 Y1.n341 0.00237961
R10570 Y1.n656 Y1.n655 0.00237961
R10571 Y1.n668 Y1.n667 0.00237961
R10572 Y1.n668 Y1.n333 0.00237961
R10573 Y1.n676 Y1.n675 0.00237961
R10574 Y1.n676 Y1.n331 0.00237961
R10575 Y1.n680 Y1.n331 0.00237961
R10576 Y1.n688 Y1.n328 0.00237961
R10577 Y1.n688 Y1.n329 0.00237961
R10578 Y1.n697 Y1.n324 0.00237961
R10579 Y1.n697 Y1.n323 0.00237961
R10580 Y1.n711 Y1.n318 0.00237961
R10581 Y1.n432 Y1.n423 0.00237961
R10582 Y1.n961 Y1.n960 0.00237961
R10583 Y1.n1022 Y1.n165 0.00237961
R10584 Y1.n1022 Y1.n1021 0.00237961
R10585 Y1.n1042 Y1.n1039 0.00237961
R10586 Y1.n143 Y1.n140 0.00237961
R10587 Y1.n1123 Y1.n114 0.00237961
R10588 Y1.n1123 Y1.n1122 0.00237961
R10589 Y1.n755 Y1.n751 0.00237961
R10590 Y1.n755 Y1.n754 0.00237961
R10591 Y1.n834 Y1.n830 0.00237961
R10592 Y1.n834 Y1.n833 0.00237961
R10593 Y1.n536 Y1.n535 0.00235952
R10594 Y1.n558 Y1.n375 0.00235952
R10595 Y1.n435 Y1.n419 0.00235749
R10596 Y1.n443 Y1.n415 0.00235749
R10597 Y1.n455 Y1.n412 0.00235749
R10598 Y1.n463 Y1.n408 0.00235749
R10599 Y1.n471 Y1.n403 0.00235749
R10600 Y1.n498 Y1.n497 0.00235749
R10601 Y1.n529 Y1.n385 0.00235749
R10602 Y1.n538 Y1.n537 0.00235749
R10603 Y1.n550 Y1.n378 0.00235749
R10604 Y1.n571 Y1.n368 0.00235749
R10605 Y1.n580 Y1.n365 0.00235749
R10606 Y1.n615 Y1.n614 0.00235749
R10607 Y1.n625 Y1.n624 0.00235749
R10608 Y1.n634 Y1.n347 0.00235749
R10609 Y1.n646 Y1.n342 0.00235749
R10610 Y1.n655 Y1.n654 0.00235749
R10611 Y1.n667 Y1.n335 0.00235749
R10612 Y1.n700 Y1.n323 0.00235749
R10613 Y1.n987 Y1.n986 0.00235749
R10614 Y1.n1093 Y1.n1092 0.00235749
R10615 Y1.n604 Y1.n603 0.00233333
R10616 Y1.n503 Y1.n498 0.00231327
R10617 Y1.n642 Y1.n344 0.00231327
R10618 Y1.n437 Y1.n436 0.00230714
R10619 Y1.n702 Y1.n322 0.00230714
R10620 Y1.n710 Y1.n703 0.00230714
R10621 Y1.n1218 Y1.n1217 0.00229115
R10622 Y1.n1307 Y1.n1306 0.00229115
R10623 Y1.n521 Y1.n388 0.00229115
R10624 Y1.n624 Y1.n351 0.00229115
R10625 Y1.n438 Y1.n416 0.00228095
R10626 Y1.n453 Y1.n409 0.00228095
R10627 Y1.n685 Y1.n684 0.00225476
R10628 Y1.n620 Y1.n615 0.00224693
R10629 Y1.n969 Y1.n968 0.00222973
R10630 Y1.n1085 Y1.n1084 0.00222973
R10631 Y1.n728 Y1.n236 0.00222973
R10632 Y1.n805 Y1.n804 0.00222973
R10633 Y1.n525 Y1.n387 0.00222482
R10634 Y1.n638 Y1.n345 0.00222482
R10635 Y1.n507 Y1.n394 0.0022027
R10636 Y1.n554 Y1.n553 0.00220238
R10637 Y1.n588 Y1.n586 0.00220238
R10638 Y1.n568 Y1.n567 0.00217619
R10639 Y1.n569 Y1.n366 0.00217619
R10640 Y1.n466 Y1.n405 0.00215848
R10641 Y1.n675 Y1.n672 0.00215848
R10642 Y1.n1242 Y1.n60 0.00213636
R10643 Y1.n1290 Y1.n1286 0.00213636
R10644 Y1.n488 Y1.n398 0.00213636
R10645 Y1.n654 Y1.n339 0.00213636
R10646 Y1.n1027 Y1.n157 0.00211425
R10647 Y1.n1138 Y1.n104 0.00211425
R10648 Y1.n772 Y1.n297 0.00211425
R10649 Y1.n850 Y1.n279 0.00211425
R10650 Y1.n721 Y1.n720 0.00209762
R10651 Y1.n452 Y1.n451 0.00209762
R10652 Y1.n584 Y1.n583 0.00209214
R10653 Y1.n988 Y1.n181 0.00209214
R10654 Y1.n125 Y1.n124 0.00209214
R10655 Y1.n736 Y1.n305 0.00209214
R10656 Y1.n816 Y1.n812 0.00209214
R10657 Y1.n686 Y1.n325 0.00207143
R10658 Y1.n537 Y1.n382 0.00207002
R10659 Y1.n557 Y1.n556 0.00207002
R10660 Y1.n605 Y1.n355 0.00204791
R10661 Y1.n435 Y1.n417 0.0020258
R10662 Y1.n701 Y1.n700 0.0020258
R10663 Y1.n711 Y1.n321 0.0020258
R10664 Y1.n541 Y1.n540 0.00201905
R10665 Y1.n983 Y1.n176 0.00201351
R10666 Y1.n1096 Y1.n1095 0.00201351
R10667 Y1.n741 Y1.n240 0.00201351
R10668 Y1.n285 Y1.n261 0.00201351
R10669 Y1.n1200 Y1.n1199 0.00200369
R10670 Y1.n1324 Y1.n35 0.00200369
R10671 Y1.n442 Y1.n439 0.00200369
R10672 Y1.n413 Y1.n410 0.00200369
R10673 Y1.n431 Y1.n429 0.00200107
R10674 Y1.n430 Y1.n193 0.00200107
R10675 Y1.n717 Y1.n317 0.00200107
R10676 Y1.n596 Y1.n356 0.00199286
R10677 Y1.n683 Y1.n328 0.00198157
R10678 Y1.n555 Y1.n376 0.00193735
R10679 Y1.n589 Y1.n362 0.00193735
R10680 Y1.n566 Y1.n368 0.00191523
R10681 Y1.n369 Y1.n367 0.00191523
R10682 Y1.n432 Y1.n420 0.00191523
R10683 Y1.n423 Y1.n422 0.00191523
R10684 Y1.n716 Y1.n319 0.00191523
R10685 Y1.n1341 Y1.n1340 0.00191523
R10686 Y1.n479 Y1.n399 0.00191429
R10687 Y1.n658 Y1.n657 0.00191429
R10688 Y1.n492 Y1.n491 0.00187101
R10689 Y1.n986 Y1.n985 0.00185493
R10690 Y1.n1093 Y1.n122 0.00185493
R10691 Y1.n1264 Y1.n1263 0.00184889
R10692 Y1.n1271 Y1.n46 0.00184889
R10693 Y1.n450 Y1.n412 0.00184889
R10694 Y1.n650 Y1.n649 0.00184889
R10695 Y1.n962 Y1.n194 0.00184889
R10696 Y1.n1060 Y1.n1059 0.00184889
R10697 Y1.n1066 Y1.n144 0.00184889
R10698 Y1.n1169 Y1.n94 0.00184889
R10699 Y1.n722 Y1.n309 0.00184889
R10700 Y1.n784 Y1.n292 0.00184889
R10701 Y1.n799 Y1.n795 0.00184889
R10702 Y1.n1343 Y1.n27 0.00184889
R10703 Y1.n629 Y1.n346 0.00183571
R10704 Y1.n329 Y1.n326 0.00182678
R10705 Y1.n511 Y1.n510 0.00180952
R10706 Y1.n1230 Y1.n66 0.0017973
R10707 Y1.n1297 Y1.n10 0.0017973
R10708 Y1.n500 Y1.n391 0.0017973
R10709 Y1.n633 Y1.n223 0.0017973
R10710 Y1.n960 Y1.n190 0.0017897
R10711 Y1.n141 Y1.n140 0.0017897
R10712 Y1.n533 Y1.n532 0.00178256
R10713 Y1.n539 Y1.n380 0.00178256
R10714 Y1.n609 Y1.n608 0.00178256
R10715 Y1.n597 Y1.n357 0.00176044
R10716 Y1.n1149 Y1.n1148 0.00175714
R10717 Y1.n512 Y1.n389 0.00173095
R10718 Y1.n628 Y1.n627 0.00173095
R10719 Y1.n459 Y1.n458 0.00171622
R10720 Y1.n1040 Y1.n1039 0.00171347
R10721 Y1.n1188 Y1.n1187 0.0016941
R10722 Y1.n1335 Y1.n1331 0.0016941
R10723 Y1.n480 Y1.n400 0.0016941
R10724 Y1.n656 Y1.n337 0.0016941
R10725 Y1.n682 Y1.n681 0.0016941
R10726 Y1.n660 Y1.n659 0.00165238
R10727 Y1.n565 Y1.n371 0.00162776
R10728 Y1.n575 Y1.n574 0.00162776
R10729 Y1.n630 Y1.n347 0.00162776
R10730 Y1.n713 Y1.n315 0.00162776
R10731 Y1.n478 Y1.n477 0.00162619
R10732 Y1.n509 Y1.n392 0.00160565
R10733 Y1.n965 Y1.n188 0.00158354
R10734 Y1.n1087 Y1.n1086 0.00158354
R10735 Y1.n729 Y1.n308 0.00158354
R10736 Y1.n803 Y1.n802 0.00158354
R10737 Y1.n1257 Y1.n51 0.00156143
R10738 Y1.n1278 Y1.n45 0.00156143
R10739 Y1.n449 Y1.n448 0.00156143
R10740 Y1.n692 Y1.n691 0.00156143
R10741 Y1.n1044 Y1.n1043 0.00156143
R10742 Y1.n1147 Y1.n1146 0.00156143
R10743 Y1.n781 Y1.n780 0.00156143
R10744 Y1.n858 Y1.n857 0.00156143
R10745 Y1.n543 Y1.n542 0.00154762
R10746 Y1.n595 Y1.n594 0.00154762
R10747 Y1.n513 Y1.n390 0.00153931
R10748 Y1.n626 Y1.n349 0.00153931
R10749 Y1.n545 Y1.n544 0.00149509
R10750 Y1.n1145 Y1.n1144 0.00149509
R10751 Y1.n598 Y1.n358 0.00147297
R10752 Y1.n661 Y1.n335 0.00147297
R10753 Y1.n446 Y1.n414 0.00146905
R10754 Y1.n694 Y1.n693 0.00146905
R10755 Y1.n476 Y1.n401 0.00145086
R10756 Y1.n1210 Y1.n74 0.00140663
R10757 Y1.n1317 Y1.n36 0.00140663
R10758 Y1.n481 Y1.n401 0.00140663
R10759 Y1.n662 Y1.n661 0.00140663
R10760 Y1.n577 Y1.n576 0.00139048
R10761 Y1.n544 Y1.n378 0.00138452
R10762 Y1.n593 Y1.n358 0.00138452
R10763 Y1.n438 Y1.n437 0.00136429
R10764 Y1.n554 Y1.n375 0.00136429
R10765 Y1.n560 Y1.n370 0.00136429
R10766 Y1.n514 Y1.n513 0.00134029
R10767 Y1.n631 Y1.n349 0.00134029
R10768 Y1.n586 Y1.n585 0.00133809
R10769 Y1.n703 Y1.n702 0.00133809
R10770 Y1.n448 Y1.n447 0.00131818
R10771 Y1.n692 Y1.n324 0.00131818
R10772 Y1.n1043 Y1.n1042 0.00131818
R10773 Y1.n743 Y1.n304 0.00129607
R10774 Y1.n765 Y1.n299 0.00129607
R10775 Y1.n820 Y1.n819 0.00129607
R10776 Y1.n843 Y1.n280 0.00129607
R10777 Y1.n461 Y1.n460 0.00128571
R10778 Y1.n679 Y1.n330 0.00128571
R10779 Y1.n1236 Y1.n62 0.00125184
R10780 Y1.n1294 Y1.n1293 0.00125184
R10781 Y1.n514 Y1.n392 0.00125184
R10782 Y1.n575 Y1.n365 0.00125184
R10783 Y1.n631 Y1.n630 0.00125184
R10784 Y1.n439 Y1.n417 0.00122973
R10785 Y1.n556 Y1.n555 0.00122973
R10786 Y1.n374 Y1.n371 0.00122973
R10787 Y1.n584 Y1.n362 0.00120762
R10788 Y1.n701 Y1.n321 0.00120762
R10789 Y1.n534 Y1.n383 0.00120714
R10790 Y1.n611 Y1.n354 0.00120714
R10791 Y1.n481 Y1.n480 0.0011855
R10792 Y1.n662 Y1.n337 0.0011855
R10793 Y1.n459 Y1.n408 0.00116339
R10794 Y1.n681 Y1.n680 0.00116339
R10795 Y1.n977 Y1.n186 0.00114865
R10796 Y1.n1081 Y1.n1077 0.00114865
R10797 Y1.n733 Y1.n732 0.00114865
R10798 Y1.n807 Y1.n259 0.00114865
R10799 Y1.n651 Y1.n340 0.00112857
R10800 Y1.n598 Y1.n597 0.00111916
R10801 Y1.n494 Y1.n397 0.00110238
R10802 Y1.n1232 Y1.n1231 0.00109705
R10803 Y1.n1299 Y1.n1298 0.00109705
R10804 Y1.n533 Y1.n384 0.00109705
R10805 Y1.n545 Y1.n380 0.00109705
R10806 Y1.n610 Y1.n609 0.00109705
R10807 Y1.n1144 Y1.n1141 0.00109705
R10808 Y1.n761 Y1.n760 0.00105283
R10809 Y1.n839 Y1.n838 0.00105283
R10810 Y1.n1340 Y1.n31 0.00105283
R10811 Y1.n1267 Y1.n1266 0.00104054
R10812 Y1.n564 Y1.n214 0.00104054
R10813 Y1.n450 Y1.n449 0.00103071
R10814 Y1.n650 Y1.n341 0.00103071
R10815 Y1.n691 Y1.n326 0.00103071
R10816 Y1.n427 Y1.n420 0.00103071
R10817 Y1.n962 Y1.n961 0.00103071
R10818 Y1.n144 Y1.n143 0.00103071
R10819 Y1.n706 Y1.n319 0.00103071
R10820 Y1.n746 Y1.n745 0.00103071
R10821 Y1.n826 Y1.n825 0.00103071
R10822 Y1.n493 Y1.n492 0.0010086
R10823 Y1.n566 Y1.n565 0.000964373
R10824 Y1.n574 Y1.n367 0.000964373
R10825 Y1.n422 Y1.n421 0.000964373
R10826 Y1.n1175 Y1.n1174 0.000964373
R10827 Y1.n713 Y1.n316 0.000964373
R10828 Y1.n1212 Y1.n72 0.00094226
R10829 Y1.n1313 Y1.n1312 0.00094226
R10830 Y1.n187 Y1.n182 0.000932432
R10831 Y1.n1078 Y1.n123 0.000932432
R10832 Y1.n737 Y1.n239 0.000932432
R10833 Y1.n813 Y1.n260 0.000932432
R10834 Y1.n432 Y1.n419 0.000898034
R10835 Y1.n683 Y1.n682 0.000898034
R10836 Y1.n458 Y1.n410 0.000875921
R10837 Y1.n716 Y1.n318 0.000853808
R10838 Y1.n1156 Y1.n1155 0.000831695
R10839 Y1.n1153 Y1.n1152 0.000814286
R10840 Y1.n532 Y1.n382 0.000809582
R10841 Y1.n608 Y1.n605 0.000809582
R10842 Y1.n1246 Y1.n1244 0.000787469
R10843 Y1.n1281 Y1.n1280 0.000787469
R10844 Y1.n988 Y1.n987 0.000787469
R10845 Y1.n1092 Y1.n124 0.000787469
R10846 Y1.n1140 Y1.n105 0.000765356
R10847 Y1.n731 Y1.n306 0.000765356
R10848 Y1.n776 Y1.n296 0.000765356
R10849 Y1.n809 Y1.n808 0.000765356
R10850 Y1.n853 Y1.n273 0.000765356
R10851 Y1.n649 Y1.n339 0.000743243
R10852 Y1.n491 Y1.n488 0.00072113
R10853 Y1.n1202 Y1.n79 0.000716216
R10854 Y1.n1327 Y1.n34 0.000716216
R10855 Y1.n457 Y1.n200 0.000716216
R10856 Y1.n327 Y1.n229 0.000716216
R10857 Y1.n502 Y1.n394 0.000676904
R10858 Y1.n1194 Y1.n1193 0.000654791
R10859 Y1.n1325 Y1.n33 0.000654791
R10860 Y1.n639 Y1.n638 0.000654791
R10861 Y1.n619 Y1.n351 0.000588452
R10862 Y1.n522 Y1.n521 0.000566339
R10863 Y1.n95 Y1.n88 0.000522113
R10864 Y1.n472 Y1.n471 0.000522113
R10865 Y2.n3 Y2.n0 15.1827
R10866 Y2.n2 Y2.n1 15.0005
R10867 Y2 Y2.n3 9.43874
R10868 Y2.n240 Y2.n239 2.2505
R10869 Y2.n241 Y2.n228 2.2505
R10870 Y2.n844 Y2.n220 2.2505
R10871 Y2.n840 Y2.n212 2.2505
R10872 Y2.n942 Y2.n941 2.2505
R10873 Y2.n948 Y2.n947 2.2505
R10874 Y2.n970 Y2.n173 2.2505
R10875 Y2.n171 Y2.n170 2.2505
R10876 Y2.n1000 Y2.n999 2.2505
R10877 Y2.n1038 Y2.n1037 2.2505
R10878 Y2.n1050 Y2.n1049 2.2505
R10879 Y2.n1045 Y2.n135 2.2505
R10880 Y2.n1043 Y2.n126 2.2505
R10881 Y2.n1142 Y2.n1141 2.2505
R10882 Y2.n1148 Y2.n1147 2.2505
R10883 Y2.n838 Y2.n240 2.2505
R10884 Y2.n847 Y2.n241 2.2505
R10885 Y2.n844 Y2.n839 2.2505
R10886 Y2.n841 Y2.n840 2.2505
R10887 Y2.n943 Y2.n942 2.2505
R10888 Y2.n947 Y2.n946 2.2505
R10889 Y2.n173 Y2.n172 2.2505
R10890 Y2.n997 Y2.n171 2.2505
R10891 Y2.n999 Y2.n998 2.2505
R10892 Y2.n1039 Y2.n1038 2.2505
R10893 Y2.n1049 Y2.n1048 2.2505
R10894 Y2.n1046 Y2.n1045 2.2505
R10895 Y2.n1043 Y2.n1042 2.2505
R10896 Y2.n1143 Y2.n1142 2.2505
R10897 Y2.n1147 Y2.n1146 2.2505
R10898 Y2.n41 Y2.n29 2.2505
R10899 Y2.n504 Y2.n32 2.2505
R10900 Y2.n658 Y2.n499 2.2505
R10901 Y2.n662 Y2.n496 2.2505
R10902 Y2.n664 Y2.n494 2.2505
R10903 Y2.n668 Y2.n491 2.2505
R10904 Y2.n670 Y2.n489 2.2505
R10905 Y2.n522 Y2.n487 2.2505
R10906 Y2.n675 Y2.n485 2.2505
R10907 Y2.n584 Y2.n482 2.2505
R10908 Y2.n681 Y2.n480 2.2505
R10909 Y2.n560 Y2.n477 2.2505
R10910 Y2.n687 Y2.n475 2.2505
R10911 Y2.n538 Y2.n470 2.2505
R10912 Y2.n469 Y2.n468 2.2505
R10913 Y2.n1346 Y2.n29 2.2505
R10914 Y2.n32 Y2.n31 2.2505
R10915 Y2.n659 Y2.n658 2.2505
R10916 Y2.n662 Y2.n661 2.2505
R10917 Y2.n665 Y2.n664 2.2505
R10918 Y2.n668 Y2.n667 2.2505
R10919 Y2.n671 Y2.n670 2.2505
R10920 Y2.n672 Y2.n487 2.2505
R10921 Y2.n675 Y2.n483 2.2505
R10922 Y2.n678 Y2.n482 2.2505
R10923 Y2.n681 Y2.n478 2.2505
R10924 Y2.n684 Y2.n477 2.2505
R10925 Y2.n687 Y2.n473 2.2505
R10926 Y2.n690 Y2.n470 2.2505
R10927 Y2.n472 Y2.n469 2.2505
R10928 Y2.n705 Y2.n454 2.2505
R10929 Y2.n706 Y2.n453 2.2505
R10930 Y2.n452 Y2.n436 2.2505
R10931 Y2.n719 Y2.n435 2.2505
R10932 Y2.n720 Y2.n434 2.2505
R10933 Y2.n433 Y2.n418 2.2505
R10934 Y2.n731 Y2.n417 2.2505
R10935 Y2.n732 Y2.n416 2.2505
R10936 Y2.n415 Y2.n402 2.2505
R10937 Y2.n414 Y2.n413 2.2505
R10938 Y2.n403 Y2.n383 2.2505
R10939 Y2.n745 Y2.n382 2.2505
R10940 Y2.n746 Y2.n381 2.2505
R10941 Y2.n380 Y2.n374 2.2505
R10942 Y2.n379 Y2.n378 2.2505
R10943 Y2.n377 Y2.n376 2.2505
R10944 Y2.n375 Y2.n352 2.2505
R10945 Y2.n769 Y2.n351 2.2505
R10946 Y2.n770 Y2.n350 2.2505
R10947 Y2.n349 Y2.n336 2.2505
R10948 Y2.n783 Y2.n335 2.2505
R10949 Y2.n784 Y2.n334 2.2505
R10950 Y2.n333 Y2.n318 2.2505
R10951 Y2.n795 Y2.n317 2.2505
R10952 Y2.n796 Y2.n316 2.2505
R10953 Y2.n315 Y2.n302 2.2505
R10954 Y2.n314 Y2.n313 2.2505
R10955 Y2.n303 Y2.n283 2.2505
R10956 Y2.n809 Y2.n282 2.2505
R10957 Y2.n810 Y2.n281 2.2505
R10958 Y2.n280 Y2.n275 2.2505
R10959 Y2.n279 Y2.n278 2.2505
R10960 Y2.n277 Y2.n276 2.2505
R10961 Y2.n243 Y2.n242 2.2505
R10962 Y2.n262 Y2.n243 2.2505
R10963 Y2.n277 Y2.n267 2.2505
R10964 Y2.n278 Y2.n268 2.2505
R10965 Y2.n275 Y2.n270 2.2505
R10966 Y2.n811 Y2.n810 2.2505
R10967 Y2.n809 Y2.n808 2.2505
R10968 Y2.n304 Y2.n283 2.2505
R10969 Y2.n313 Y2.n312 2.2505
R10970 Y2.n302 Y2.n300 2.2505
R10971 Y2.n797 Y2.n796 2.2505
R10972 Y2.n795 Y2.n794 2.2505
R10973 Y2.n330 Y2.n318 2.2505
R10974 Y2.n785 Y2.n784 2.2505
R10975 Y2.n783 Y2.n782 2.2505
R10976 Y2.n345 Y2.n336 2.2505
R10977 Y2.n771 Y2.n770 2.2505
R10978 Y2.n769 Y2.n768 2.2505
R10979 Y2.n363 Y2.n352 2.2505
R10980 Y2.n377 Y2.n367 2.2505
R10981 Y2.n378 Y2.n368 2.2505
R10982 Y2.n374 Y2.n370 2.2505
R10983 Y2.n747 Y2.n746 2.2505
R10984 Y2.n745 Y2.n744 2.2505
R10985 Y2.n404 Y2.n383 2.2505
R10986 Y2.n413 Y2.n412 2.2505
R10987 Y2.n402 Y2.n400 2.2505
R10988 Y2.n733 Y2.n732 2.2505
R10989 Y2.n731 Y2.n730 2.2505
R10990 Y2.n430 Y2.n418 2.2505
R10991 Y2.n721 Y2.n720 2.2505
R10992 Y2.n719 Y2.n718 2.2505
R10993 Y2.n448 Y2.n436 2.2505
R10994 Y2.n707 Y2.n706 2.2505
R10995 Y2.n705 Y2.n704 2.2505
R10996 Y2.n1163 Y2.n95 2.2505
R10997 Y2.n1176 Y2.n1175 2.2505
R10998 Y2.n100 Y2.n92 2.2505
R10999 Y2.n1186 Y2.n1185 2.2505
R11000 Y2.n93 Y2.n89 2.2505
R11001 Y2.n1181 Y2.n87 2.2505
R11002 Y2.n1180 Y2.n85 2.2505
R11003 Y2.n1200 Y2.n79 2.2505
R11004 Y2.n1216 Y2.n1215 2.2505
R11005 Y2.n1208 Y2.n77 2.2505
R11006 Y2.n1221 Y2.n1220 2.2505
R11007 Y2.n1224 Y2.n69 2.2505
R11008 Y2.n1237 Y2.n1236 2.2505
R11009 Y2.n71 Y2.n67 2.2505
R11010 Y2.n1242 Y2.n1241 2.2505
R11011 Y2.n1251 Y2.n6 2.2505
R11012 Y2.n1374 Y2.n7 2.2505
R11013 Y2.n1373 Y2.n8 2.2505
R11014 Y2.n1372 Y2.n9 2.2505
R11015 Y2.n1269 Y2.n10 2.2505
R11016 Y2.n1368 Y2.n12 2.2505
R11017 Y2.n1367 Y2.n13 2.2505
R11018 Y2.n1366 Y2.n14 2.2505
R11019 Y2.n1286 Y2.n15 2.2505
R11020 Y2.n1362 Y2.n17 2.2505
R11021 Y2.n1361 Y2.n18 2.2505
R11022 Y2.n1360 Y2.n19 2.2505
R11023 Y2.n50 Y2.n20 2.2505
R11024 Y2.n1356 Y2.n22 2.2505
R11025 Y2.n1355 Y2.n23 2.2505
R11026 Y2.n1354 Y2.n24 2.2505
R11027 Y2.n1325 Y2.n25 2.2505
R11028 Y2.n1350 Y2.n27 2.2505
R11029 Y2.n1349 Y2.n28 2.2505
R11030 Y2.n1349 Y2.n26 2.2505
R11031 Y2.n1351 Y2.n1350 2.2505
R11032 Y2.n1352 Y2.n25 2.2505
R11033 Y2.n1354 Y2.n1353 2.2505
R11034 Y2.n1355 Y2.n21 2.2505
R11035 Y2.n1357 Y2.n1356 2.2505
R11036 Y2.n1358 Y2.n20 2.2505
R11037 Y2.n1360 Y2.n1359 2.2505
R11038 Y2.n1361 Y2.n16 2.2505
R11039 Y2.n1363 Y2.n1362 2.2505
R11040 Y2.n1364 Y2.n15 2.2505
R11041 Y2.n1366 Y2.n1365 2.2505
R11042 Y2.n1367 Y2.n11 2.2505
R11043 Y2.n1369 Y2.n1368 2.2505
R11044 Y2.n1370 Y2.n10 2.2505
R11045 Y2.n1372 Y2.n1371 2.2505
R11046 Y2.n1373 Y2.n5 2.2505
R11047 Y2.n1375 Y2.n1374 2.2505
R11048 Y2.n6 Y2.n4 2.2505
R11049 Y2.n1241 Y2.n1240 2.2505
R11050 Y2.n1239 Y2.n67 2.2505
R11051 Y2.n1238 Y2.n1237 2.2505
R11052 Y2.n69 Y2.n68 2.2505
R11053 Y2.n1220 Y2.n1219 2.2505
R11054 Y2.n1218 Y2.n77 2.2505
R11055 Y2.n1217 Y2.n1216 2.2505
R11056 Y2.n79 Y2.n78 2.2505
R11057 Y2.n1180 Y2.n1179 2.2505
R11058 Y2.n1182 Y2.n1181 2.2505
R11059 Y2.n1183 Y2.n93 2.2505
R11060 Y2.n1185 Y2.n1184 2.2505
R11061 Y2.n1178 Y2.n92 2.2505
R11062 Y2.n1177 Y2.n1176 2.2505
R11063 Y2.n95 Y2.n94 2.2505
R11064 Y2.n1150 Y2.n1149 2.2005
R11065 Y2.n1123 Y2.n113 2.2005
R11066 Y2.n1127 Y2.n1118 2.2005
R11067 Y2.n1116 Y2.n1114 2.2005
R11068 Y2.n1134 Y2.n119 2.2005
R11069 Y2.n1140 Y2.n1139 2.2005
R11070 Y2.n1109 Y2.n118 2.2005
R11071 Y2.n1100 Y2.n123 2.2005
R11072 Y2.n1103 Y2.n1102 2.2005
R11073 Y2.n1099 Y2.n1098 2.2005
R11074 Y2.n1092 Y2.n1091 2.2005
R11075 Y2.n1090 Y2.n1089 2.2005
R11076 Y2.n1083 Y2.n1082 2.2005
R11077 Y2.n1081 Y2.n1080 2.2005
R11078 Y2.n1075 Y2.n1074 2.2005
R11079 Y2.n1073 Y2.n1072 2.2005
R11080 Y2.n1067 Y2.n1066 2.2005
R11081 Y2.n1065 Y2.n1064 2.2005
R11082 Y2.n1058 Y2.n144 2.2005
R11083 Y2.n1052 Y2.n1051 2.2005
R11084 Y2.n150 Y2.n149 2.2005
R11085 Y2.n1030 Y2.n157 2.2005
R11086 Y2.n1036 Y2.n1035 2.2005
R11087 Y2.n1024 Y2.n155 2.2005
R11088 Y2.n1018 Y2.n1017 2.2005
R11089 Y2.n1015 Y2.n1014 2.2005
R11090 Y2.n1010 Y2.n164 2.2005
R11091 Y2.n1001 Y2.n167 2.2005
R11092 Y2.n1003 Y2.n1002 2.2005
R11093 Y2.n987 Y2.n175 2.2005
R11094 Y2.n993 Y2.n992 2.2005
R11095 Y2.n980 Y2.n174 2.2005
R11096 Y2.n971 Y2.n179 2.2005
R11097 Y2.n973 Y2.n972 2.2005
R11098 Y2.n969 Y2.n968 2.2005
R11099 Y2.n962 Y2.n182 2.2005
R11100 Y2.n194 Y2.n186 2.2005
R11101 Y2.n955 Y2.n189 2.2005
R11102 Y2.n950 Y2.n949 2.2005
R11103 Y2.n933 Y2.n192 2.2005
R11104 Y2.n203 Y2.n201 2.2005
R11105 Y2.n940 Y2.n939 2.2005
R11106 Y2.n926 Y2.n199 2.2005
R11107 Y2.n920 Y2.n919 2.2005
R11108 Y2.n918 Y2.n917 2.2005
R11109 Y2.n912 Y2.n911 2.2005
R11110 Y2.n910 Y2.n909 2.2005
R11111 Y2.n905 Y2.n904 2.2005
R11112 Y2.n903 Y2.n902 2.2005
R11113 Y2.n896 Y2.n895 2.2005
R11114 Y2.n894 Y2.n893 2.2005
R11115 Y2.n886 Y2.n885 2.2005
R11116 Y2.n884 Y2.n883 2.2005
R11117 Y2.n877 Y2.n876 2.2005
R11118 Y2.n875 Y2.n874 2.2005
R11119 Y2.n869 Y2.n868 2.2005
R11120 Y2.n867 Y2.n866 2.2005
R11121 Y2.n860 Y2.n232 2.2005
R11122 Y2.n851 Y2.n236 2.2005
R11123 Y2.n853 Y2.n852 2.2005
R11124 Y2.n253 Y2.n244 2.2005
R11125 Y2.n43 Y2.n42 2.2005
R11126 Y2.n463 Y2.n457 2.2005
R11127 Y2.n466 Y2.n464 2.2005
R11128 Y2.n695 Y2.n694 2.2005
R11129 Y2.n467 Y2.n465 2.2005
R11130 Y2.n541 Y2.n540 2.2005
R11131 Y2.n543 Y2.n542 2.2005
R11132 Y2.n545 Y2.n544 2.2005
R11133 Y2.n547 Y2.n546 2.2005
R11134 Y2.n549 Y2.n548 2.2005
R11135 Y2.n551 Y2.n550 2.2005
R11136 Y2.n553 Y2.n552 2.2005
R11137 Y2.n555 Y2.n554 2.2005
R11138 Y2.n558 Y2.n557 2.2005
R11139 Y2.n559 Y2.n533 2.2005
R11140 Y2.n563 Y2.n562 2.2005
R11141 Y2.n561 Y2.n531 2.2005
R11142 Y2.n569 Y2.n568 2.2005
R11143 Y2.n570 Y2.n530 2.2005
R11144 Y2.n572 Y2.n571 2.2005
R11145 Y2.n575 Y2.n574 2.2005
R11146 Y2.n577 Y2.n576 2.2005
R11147 Y2.n528 Y2.n527 2.2005
R11148 Y2.n583 Y2.n582 2.2005
R11149 Y2.n585 Y2.n526 2.2005
R11150 Y2.n587 Y2.n586 2.2005
R11151 Y2.n589 Y2.n588 2.2005
R11152 Y2.n591 Y2.n590 2.2005
R11153 Y2.n593 Y2.n592 2.2005
R11154 Y2.n596 Y2.n595 2.2005
R11155 Y2.n594 Y2.n523 2.2005
R11156 Y2.n602 Y2.n601 2.2005
R11157 Y2.n604 Y2.n603 2.2005
R11158 Y2.n606 Y2.n605 2.2005
R11159 Y2.n608 Y2.n607 2.2005
R11160 Y2.n610 Y2.n609 2.2005
R11161 Y2.n612 Y2.n611 2.2005
R11162 Y2.n614 Y2.n613 2.2005
R11163 Y2.n616 Y2.n615 2.2005
R11164 Y2.n518 Y2.n517 2.2005
R11165 Y2.n622 Y2.n621 2.2005
R11166 Y2.n624 Y2.n516 2.2005
R11167 Y2.n626 Y2.n625 2.2005
R11168 Y2.n629 Y2.n628 2.2005
R11169 Y2.n630 Y2.n515 2.2005
R11170 Y2.n632 Y2.n631 2.2005
R11171 Y2.n635 Y2.n634 2.2005
R11172 Y2.n633 Y2.n513 2.2005
R11173 Y2.n640 Y2.n512 2.2005
R11174 Y2.n643 Y2.n642 2.2005
R11175 Y2.n645 Y2.n511 2.2005
R11176 Y2.n647 Y2.n646 2.2005
R11177 Y2.n649 Y2.n648 2.2005
R11178 Y2.n502 Y2.n500 2.2005
R11179 Y2.n655 Y2.n654 2.2005
R11180 Y2.n509 Y2.n501 2.2005
R11181 Y2.n508 Y2.n507 2.2005
R11182 Y2.n506 Y2.n505 2.2005
R11183 Y2.n35 Y2.n33 2.2005
R11184 Y2.n1342 Y2.n1341 2.2005
R11185 Y2.n36 Y2.n34 2.2005
R11186 Y2.n829 Y2.n245 2.2005
R11187 Y2.n827 Y2.n263 2.2005
R11188 Y2.n266 Y2.n264 2.2005
R11189 Y2.n822 Y2.n821 2.2005
R11190 Y2.n820 Y2.n819 2.2005
R11191 Y2.n818 Y2.n817 2.2005
R11192 Y2.n816 Y2.n815 2.2005
R11193 Y2.n813 Y2.n812 2.2005
R11194 Y2.n290 Y2.n274 2.2005
R11195 Y2.n291 Y2.n284 2.2005
R11196 Y2.n807 Y2.n806 2.2005
R11197 Y2.n287 Y2.n285 2.2005
R11198 Y2.n306 Y2.n305 2.2005
R11199 Y2.n308 Y2.n307 2.2005
R11200 Y2.n311 Y2.n310 2.2005
R11201 Y2.n309 Y2.n298 2.2005
R11202 Y2.n800 Y2.n799 2.2005
R11203 Y2.n798 Y2.n299 2.2005
R11204 Y2.n323 Y2.n301 2.2005
R11205 Y2.n325 Y2.n319 2.2005
R11206 Y2.n793 Y2.n792 2.2005
R11207 Y2.n327 Y2.n320 2.2005
R11208 Y2.n331 Y2.n328 2.2005
R11209 Y2.n787 Y2.n786 2.2005
R11210 Y2.n332 Y2.n329 2.2005
R11211 Y2.n340 Y2.n337 2.2005
R11212 Y2.n781 Y2.n780 2.2005
R11213 Y2.n342 Y2.n338 2.2005
R11214 Y2.n775 Y2.n346 2.2005
R11215 Y2.n773 Y2.n772 2.2005
R11216 Y2.n356 Y2.n348 2.2005
R11217 Y2.n357 Y2.n353 2.2005
R11218 Y2.n767 Y2.n766 2.2005
R11219 Y2.n358 Y2.n354 2.2005
R11220 Y2.n364 Y2.n362 2.2005
R11221 Y2.n760 Y2.n365 2.2005
R11222 Y2.n758 Y2.n757 2.2005
R11223 Y2.n756 Y2.n755 2.2005
R11224 Y2.n754 Y2.n753 2.2005
R11225 Y2.n752 Y2.n751 2.2005
R11226 Y2.n749 Y2.n748 2.2005
R11227 Y2.n390 Y2.n373 2.2005
R11228 Y2.n391 Y2.n384 2.2005
R11229 Y2.n743 Y2.n742 2.2005
R11230 Y2.n387 Y2.n385 2.2005
R11231 Y2.n406 Y2.n405 2.2005
R11232 Y2.n408 Y2.n407 2.2005
R11233 Y2.n411 Y2.n410 2.2005
R11234 Y2.n409 Y2.n398 2.2005
R11235 Y2.n736 Y2.n735 2.2005
R11236 Y2.n734 Y2.n399 2.2005
R11237 Y2.n423 Y2.n401 2.2005
R11238 Y2.n425 Y2.n419 2.2005
R11239 Y2.n729 Y2.n728 2.2005
R11240 Y2.n427 Y2.n420 2.2005
R11241 Y2.n431 Y2.n428 2.2005
R11242 Y2.n723 Y2.n722 2.2005
R11243 Y2.n432 Y2.n429 2.2005
R11244 Y2.n441 Y2.n437 2.2005
R11245 Y2.n717 Y2.n716 2.2005
R11246 Y2.n440 Y2.n438 2.2005
R11247 Y2.n710 Y2.n449 2.2005
R11248 Y2.n709 Y2.n708 2.2005
R11249 Y2.n459 Y2.n451 2.2005
R11250 Y2.n460 Y2.n456 2.2005
R11251 Y2.n1162 Y2.n1161 2.2005
R11252 Y2.n1165 Y2.n1164 2.2005
R11253 Y2.n98 Y2.n96 2.2005
R11254 Y2.n1174 Y2.n1173 2.2005
R11255 Y2.n103 Y2.n97 2.2005
R11256 Y2.n102 Y2.n101 2.2005
R11257 Y2.n99 Y2.n91 2.2005
R11258 Y2.n1188 Y2.n1187 2.2005
R11259 Y2.n1190 Y2.n1189 2.2005
R11260 Y2.n1192 Y2.n1191 2.2005
R11261 Y2.n1194 Y2.n1193 2.2005
R11262 Y2.n1196 Y2.n1195 2.2005
R11263 Y2.n1198 Y2.n1197 2.2005
R11264 Y2.n1199 Y2.n84 2.2005
R11265 Y2.n1202 Y2.n1201 2.2005
R11266 Y2.n82 Y2.n80 2.2005
R11267 Y2.n1214 Y2.n1213 2.2005
R11268 Y2.n1212 Y2.n81 2.2005
R11269 Y2.n1210 Y2.n1209 2.2005
R11270 Y2.n1207 Y2.n76 2.2005
R11271 Y2.n1222 Y2.n75 2.2005
R11272 Y2.n1226 Y2.n1225 2.2005
R11273 Y2.n1223 Y2.n73 2.2005
R11274 Y2.n1231 Y2.n70 2.2005
R11275 Y2.n1235 Y2.n1234 2.2005
R11276 Y2.n1232 Y2.n72 2.2005
R11277 Y2.n66 Y2.n65 2.2005
R11278 Y2.n1244 Y2.n1243 2.2005
R11279 Y2.n63 Y2.n62 2.2005
R11280 Y2.n1250 Y2.n1249 2.2005
R11281 Y2.n1252 Y2.n61 2.2005
R11282 Y2.n1254 Y2.n1253 2.2005
R11283 Y2.n1256 Y2.n1255 2.2005
R11284 Y2.n1258 Y2.n1257 2.2005
R11285 Y2.n1260 Y2.n1259 2.2005
R11286 Y2.n1262 Y2.n1261 2.2005
R11287 Y2.n59 Y2.n58 2.2005
R11288 Y2.n1268 Y2.n1267 2.2005
R11289 Y2.n1270 Y2.n57 2.2005
R11290 Y2.n1272 Y2.n1271 2.2005
R11291 Y2.n1275 Y2.n1274 2.2005
R11292 Y2.n1277 Y2.n1276 2.2005
R11293 Y2.n1279 Y2.n1278 2.2005
R11294 Y2.n55 Y2.n54 2.2005
R11295 Y2.n1285 Y2.n1284 2.2005
R11296 Y2.n1287 Y2.n53 2.2005
R11297 Y2.n1289 Y2.n1288 2.2005
R11298 Y2.n1292 Y2.n1291 2.2005
R11299 Y2.n1294 Y2.n1293 2.2005
R11300 Y2.n1297 Y2.n1296 2.2005
R11301 Y2.n1295 Y2.n51 2.2005
R11302 Y2.n1304 Y2.n1303 2.2005
R11303 Y2.n1306 Y2.n1305 2.2005
R11304 Y2.n1308 Y2.n1307 2.2005
R11305 Y2.n1310 Y2.n1309 2.2005
R11306 Y2.n1312 Y2.n1311 2.2005
R11307 Y2.n1314 Y2.n1313 2.2005
R11308 Y2.n1316 Y2.n1315 2.2005
R11309 Y2.n1318 Y2.n1317 2.2005
R11310 Y2.n46 Y2.n45 2.2005
R11311 Y2.n1324 Y2.n1323 2.2005
R11312 Y2.n1326 Y2.n44 2.2005
R11313 Y2.n1328 Y2.n1327 2.2005
R11314 Y2.n1331 Y2.n1330 2.2005
R11315 Y2.n1333 Y2.n1332 2.2005
R11316 Y2.n850 Y2.n849 1.8005
R11317 Y2.n845 Y2.n224 1.8005
R11318 Y2.n843 Y2.n216 1.8005
R11319 Y2.n208 Y2.n198 1.8005
R11320 Y2.n200 Y2.n193 1.8005
R11321 Y2.n196 Y2.n195 1.8005
R11322 Y2.n995 Y2.n994 1.8005
R11323 Y2.n1016 Y2.n154 1.8005
R11324 Y2.n156 Y2.n151 1.8005
R11325 Y2.n152 Y2.n140 1.8005
R11326 Y2.n1044 Y2.n130 1.8005
R11327 Y2.n1101 Y2.n117 1.8005
R11328 Y2.n1117 Y2.n114 1.8005
R11329 Y2.n849 Y2.n848 1.8005
R11330 Y2.n846 Y2.n845 1.8005
R11331 Y2.n843 Y2.n842 1.8005
R11332 Y2.n198 Y2.n197 1.8005
R11333 Y2.n944 Y2.n193 1.8005
R11334 Y2.n945 Y2.n196 1.8005
R11335 Y2.n996 Y2.n995 1.8005
R11336 Y2.n154 Y2.n153 1.8005
R11337 Y2.n1040 Y2.n151 1.8005
R11338 Y2.n1047 Y2.n152 1.8005
R11339 Y2.n1044 Y2.n1041 1.8005
R11340 Y2.n117 Y2.n116 1.8005
R11341 Y2.n1144 Y2.n114 1.8005
R11342 Y2.n1344 Y2.n1343 1.8005
R11343 Y2.n657 Y2.n656 1.8005
R11344 Y2.n644 Y2.n497 1.8005
R11345 Y2.n663 Y2.n495 1.8005
R11346 Y2.n623 Y2.n492 1.8005
R11347 Y2.n669 Y2.n490 1.8005
R11348 Y2.n674 Y2.n486 1.8005
R11349 Y2.n676 Y2.n484 1.8005
R11350 Y2.n680 Y2.n481 1.8005
R11351 Y2.n682 Y2.n479 1.8005
R11352 Y2.n686 Y2.n476 1.8005
R11353 Y2.n688 Y2.n474 1.8005
R11354 Y2.n693 Y2.n692 1.8005
R11355 Y2.n1345 Y2.n1344 1.8005
R11356 Y2.n657 Y2.n498 1.8005
R11357 Y2.n660 Y2.n497 1.8005
R11358 Y2.n663 Y2.n493 1.8005
R11359 Y2.n666 Y2.n492 1.8005
R11360 Y2.n669 Y2.n488 1.8005
R11361 Y2.n674 Y2.n673 1.8005
R11362 Y2.n677 Y2.n676 1.8005
R11363 Y2.n680 Y2.n679 1.8005
R11364 Y2.n683 Y2.n682 1.8005
R11365 Y2.n686 Y2.n685 1.8005
R11366 Y2.n689 Y2.n688 1.8005
R11367 Y2.n692 Y2.n691 1.8005
R11368 Y2.n471 Y2.n455 1.8005
R11369 Y2.n703 Y2.n455 1.8005
R11370 Y2.n1348 Y2.n30 1.8005
R11371 Y2.n1348 Y2.n1347 1.8005
R11372 Y2.n837 Y2.n836 1.5005
R11373 Y2.n836 Y2.n835 1.5005
R11374 Y2.n115 Y2.n106 1.5005
R11375 Y2.n1145 Y2.n115 1.5005
R11376 Y2.n1158 Y2.n105 1.1125
R11377 Y2.n715 Y2.n714 1.10836
R11378 Y2.n446 Y2.n439 1.10443
R11379 Y2.n700 Y2.n461 1.10381
R11380 Y2.n1160 Y2.n1159 1.10372
R11381 Y2.n442 Y2.n426 1.10339
R11382 Y2.n710 Y2.n447 1.10272
R11383 Y2.n713 Y2.n440 1.10272
R11384 Y2.n445 Y2.n441 1.10272
R11385 Y2.n1165 Y2.n104 1.10263
R11386 Y2.n1168 Y2.n98 1.10263
R11387 Y2.n1340 Y2.n1339 1.1005
R11388 Y2.n697 Y2.n696 1.1005
R11389 Y2.n539 Y2.n462 1.1005
R11390 Y2.n537 Y2.n536 1.1005
R11391 Y2.n535 Y2.n534 1.1005
R11392 Y2.n556 Y2.n532 1.1005
R11393 Y2.n565 Y2.n564 1.1005
R11394 Y2.n567 Y2.n566 1.1005
R11395 Y2.n573 Y2.n529 1.1005
R11396 Y2.n579 Y2.n578 1.1005
R11397 Y2.n581 Y2.n580 1.1005
R11398 Y2.n525 Y2.n524 1.1005
R11399 Y2.n598 Y2.n597 1.1005
R11400 Y2.n601 Y2.n600 1.1005
R11401 Y2.n599 Y2.n521 1.1005
R11402 Y2.n520 Y2.n519 1.1005
R11403 Y2.n618 Y2.n617 1.1005
R11404 Y2.n620 Y2.n619 1.1005
R11405 Y2.n627 Y2.n514 1.1005
R11406 Y2.n637 Y2.n636 1.1005
R11407 Y2.n639 Y2.n638 1.1005
R11408 Y2.n641 Y2.n510 1.1005
R11409 Y2.n651 Y2.n650 1.1005
R11410 Y2.n653 Y2.n652 1.1005
R11411 Y2.n503 Y2.n37 1.1005
R11412 Y2.n698 Y2.n458 1.1005
R11413 Y2.n825 Y2.n824 1.1005
R11414 Y2.n292 Y2.n289 1.1005
R11415 Y2.n776 Y2.n343 1.1005
R11416 Y2.n761 Y2.n360 1.1005
R11417 Y2.n392 Y2.n389 1.1005
R11418 Y2.n699 Y2.n450 1.1005
R11419 Y2.n712 Y2.n711 1.1005
R11420 Y2.n444 Y2.n443 1.1005
R11421 Y2.n725 Y2.n724 1.1005
R11422 Y2.n738 Y2.n737 1.1005
R11423 Y2.n394 Y2.n393 1.1005
R11424 Y2.n366 Y2.n361 1.1005
R11425 Y2.n763 Y2.n762 1.1005
R11426 Y2.n347 Y2.n344 1.1005
R11427 Y2.n778 Y2.n777 1.1005
R11428 Y2.n789 Y2.n788 1.1005
R11429 Y2.n802 Y2.n801 1.1005
R11430 Y2.n294 Y2.n293 1.1005
R11431 Y2.n271 Y2.n265 1.1005
R11432 Y2.n826 Y2.n261 1.1005
R11433 Y2.n832 Y2.n248 1.1005
R11434 Y2.n260 Y2.n247 1.1005
R11435 Y2.n831 Y2.n830 1.1005
R11436 Y2.n834 Y2.n833 1.1005
R11437 Y2.n1150 Y2.n111 1.1005
R11438 Y2.n1122 Y2.n1121 1.1005
R11439 Y2.n1124 Y2.n1123 1.1005
R11440 Y2.n1127 Y2.n1126 1.1005
R11441 Y2.n1130 Y2.n1129 1.1005
R11442 Y2.n1133 Y2.n1113 1.1005
R11443 Y2.n1135 Y2.n1134 1.1005
R11444 Y2.n1136 Y2.n121 1.1005
R11445 Y2.n1111 Y2.n1110 1.1005
R11446 Y2.n1096 Y2.n125 1.1005
R11447 Y2.n1098 Y2.n1097 1.1005
R11448 Y2.n1095 Y2.n127 1.1005
R11449 Y2.n1087 Y2.n132 1.1005
R11450 Y2.n1089 Y2.n1088 1.1005
R11451 Y2.n1086 Y2.n131 1.1005
R11452 Y2.n1078 Y2.n137 1.1005
R11453 Y2.n1069 Y2.n141 1.1005
R11454 Y2.n1068 Y2.n1067 1.1005
R11455 Y2.n143 Y2.n142 1.1005
R11456 Y2.n1060 Y2.n1059 1.1005
R11457 Y2.n1058 Y2.n146 1.1005
R11458 Y2.n1057 Y2.n1056 1.1005
R11459 Y2.n1054 Y2.n1053 1.1005
R11460 Y2.n149 Y2.n148 1.1005
R11461 Y2.n1031 Y2.n1030 1.1005
R11462 Y2.n1034 Y2.n1033 1.1005
R11463 Y2.n1026 Y2.n1025 1.1005
R11464 Y2.n1024 Y2.n160 1.1005
R11465 Y2.n1023 Y2.n1022 1.1005
R11466 Y2.n163 Y2.n162 1.1005
R11467 Y2.n1008 Y2.n1007 1.1005
R11468 Y2.n1006 Y2.n167 1.1005
R11469 Y2.n1003 Y2.n168 1.1005
R11470 Y2.n986 Y2.n985 1.1005
R11471 Y2.n990 Y2.n177 1.1005
R11472 Y2.n992 Y2.n991 1.1005
R11473 Y2.n983 Y2.n176 1.1005
R11474 Y2.n978 Y2.n977 1.1005
R11475 Y2.n966 Y2.n184 1.1005
R11476 Y2.n968 Y2.n967 1.1005
R11477 Y2.n963 Y2.n962 1.1005
R11478 Y2.n960 Y2.n959 1.1005
R11479 Y2.n956 Y2.n187 1.1005
R11480 Y2.n955 Y2.n954 1.1005
R11481 Y2.n953 Y2.n188 1.1005
R11482 Y2.n932 Y2.n931 1.1005
R11483 Y2.n928 Y2.n927 1.1005
R11484 Y2.n926 Y2.n204 1.1005
R11485 Y2.n925 Y2.n924 1.1005
R11486 Y2.n207 Y2.n206 1.1005
R11487 Y2.n917 Y2.n916 1.1005
R11488 Y2.n915 Y2.n209 1.1005
R11489 Y2.n211 Y2.n210 1.1005
R11490 Y2.n909 Y2.n908 1.1005
R11491 Y2.n906 Y2.n905 1.1005
R11492 Y2.n901 Y2.n900 1.1005
R11493 Y2.n898 Y2.n897 1.1005
R11494 Y2.n896 Y2.n218 1.1005
R11495 Y2.n890 Y2.n219 1.1005
R11496 Y2.n888 Y2.n887 1.1005
R11497 Y2.n886 Y2.n222 1.1005
R11498 Y2.n880 Y2.n223 1.1005
R11499 Y2.n879 Y2.n225 1.1005
R11500 Y2.n878 Y2.n877 1.1005
R11501 Y2.n874 Y2.n873 1.1005
R11502 Y2.n871 Y2.n870 1.1005
R11503 Y2.n864 Y2.n234 1.1005
R11504 Y2.n866 Y2.n865 1.1005
R11505 Y2.n863 Y2.n233 1.1005
R11506 Y2.n858 Y2.n857 1.1005
R11507 Y2.n252 Y2.n251 1.1005
R11508 Y2.n254 Y2.n253 1.1005
R11509 Y2.n258 Y2.n257 1.1005
R11510 Y2.n259 Y2.n258 1.1005
R11511 Y2.n256 Y2.n247 1.1005
R11512 Y2.n255 Y2.n246 1.1005
R11513 Y2.n856 Y2.n236 1.1005
R11514 Y2.n855 Y2.n854 1.1005
R11515 Y2.n853 Y2.n237 1.1005
R11516 Y2.n250 Y2.n238 1.1005
R11517 Y2.n859 Y2.n235 1.1005
R11518 Y2.n862 Y2.n861 1.1005
R11519 Y2.n231 Y2.n230 1.1005
R11520 Y2.n872 Y2.n229 1.1005
R11521 Y2.n227 Y2.n226 1.1005
R11522 Y2.n882 Y2.n881 1.1005
R11523 Y2.n889 Y2.n221 1.1005
R11524 Y2.n892 Y2.n891 1.1005
R11525 Y2.n899 Y2.n217 1.1005
R11526 Y2.n215 Y2.n214 1.1005
R11527 Y2.n907 Y2.n213 1.1005
R11528 Y2.n914 Y2.n913 1.1005
R11529 Y2.n922 Y2.n921 1.1005
R11530 Y2.n923 Y2.n205 1.1005
R11531 Y2.n929 Y2.n202 1.1005
R11532 Y2.n933 Y2.n930 1.1005
R11533 Y2.n935 Y2.n934 1.1005
R11534 Y2.n936 Y2.n203 1.1005
R11535 Y2.n938 Y2.n937 1.1005
R11536 Y2.n191 Y2.n190 1.1005
R11537 Y2.n952 Y2.n951 1.1005
R11538 Y2.n958 Y2.n957 1.1005
R11539 Y2.n961 Y2.n185 1.1005
R11540 Y2.n964 Y2.n183 1.1005
R11541 Y2.n976 Y2.n179 1.1005
R11542 Y2.n975 Y2.n974 1.1005
R11543 Y2.n973 Y2.n180 1.1005
R11544 Y2.n965 Y2.n181 1.1005
R11545 Y2.n979 Y2.n178 1.1005
R11546 Y2.n982 Y2.n981 1.1005
R11547 Y2.n989 Y2.n988 1.1005
R11548 Y2.n984 Y2.n169 1.1005
R11549 Y2.n1005 Y2.n1004 1.1005
R11550 Y2.n1014 Y2.n1013 1.1005
R11551 Y2.n1012 Y2.n165 1.1005
R11552 Y2.n1011 Y2.n1010 1.1005
R11553 Y2.n1009 Y2.n166 1.1005
R11554 Y2.n1020 Y2.n1019 1.1005
R11555 Y2.n1021 Y2.n161 1.1005
R11556 Y2.n1027 Y2.n158 1.1005
R11557 Y2.n1032 Y2.n159 1.1005
R11558 Y2.n1029 Y2.n1028 1.1005
R11559 Y2.n1055 Y2.n147 1.1005
R11560 Y2.n1061 Y2.n145 1.1005
R11561 Y2.n1063 Y2.n1062 1.1005
R11562 Y2.n1071 Y2.n1070 1.1005
R11563 Y2.n1080 Y2.n1079 1.1005
R11564 Y2.n1077 Y2.n136 1.1005
R11565 Y2.n1076 Y2.n1075 1.1005
R11566 Y2.n139 Y2.n138 1.1005
R11567 Y2.n134 Y2.n133 1.1005
R11568 Y2.n1085 Y2.n1084 1.1005
R11569 Y2.n129 Y2.n128 1.1005
R11570 Y2.n1094 Y2.n1093 1.1005
R11571 Y2.n1103 Y2.n124 1.1005
R11572 Y2.n1109 Y2.n122 1.1005
R11573 Y2.n1108 Y2.n1107 1.1005
R11574 Y2.n1106 Y2.n123 1.1005
R11575 Y2.n1105 Y2.n1104 1.1005
R11576 Y2.n1112 Y2.n120 1.1005
R11577 Y2.n1138 Y2.n1137 1.1005
R11578 Y2.n1132 Y2.n1131 1.1005
R11579 Y2.n1128 Y2.n1115 1.1005
R11580 Y2.n1125 Y2.n1119 1.1005
R11581 Y2.n1120 Y2.n112 1.1005
R11582 Y2.n1152 Y2.n1151 1.1005
R11583 Y2.n1156 Y2.n1155 1.1005
R11584 Y2.n109 Y2.n108 1.1005
R11585 Y2.n39 Y2.n38 1.1005
R11586 Y2.n1337 Y2.n1336 1.1005
R11587 Y2.n1338 Y2.n1337 1.1005
R11588 Y2.n1155 Y2.n1154 1.1005
R11589 Y2.n1153 Y2.n109 1.1005
R11590 Y2.n1335 Y2.n1334 1.1005
R11591 Y2.n1329 Y2.n40 1.1005
R11592 Y2.n1322 Y2.n1321 1.1005
R11593 Y2.n1320 Y2.n1319 1.1005
R11594 Y2.n48 Y2.n47 1.1005
R11595 Y2.n1300 Y2.n49 1.1005
R11596 Y2.n1302 Y2.n1301 1.1005
R11597 Y2.n1299 Y2.n1298 1.1005
R11598 Y2.n1290 Y2.n52 1.1005
R11599 Y2.n1283 Y2.n1282 1.1005
R11600 Y2.n1281 Y2.n1280 1.1005
R11601 Y2.n1273 Y2.n56 1.1005
R11602 Y2.n1266 Y2.n1265 1.1005
R11603 Y2.n1264 Y2.n1263 1.1005
R11604 Y2.n1255 Y2.n60 1.1005
R11605 Y2.n1248 Y2.n1247 1.1005
R11606 Y2.n1246 Y2.n1245 1.1005
R11607 Y2.n1233 Y2.n64 1.1005
R11608 Y2.n1230 Y2.n1229 1.1005
R11609 Y2.n1228 Y2.n1227 1.1005
R11610 Y2.n1211 Y2.n74 1.1005
R11611 Y2.n1206 Y2.n1205 1.1005
R11612 Y2.n1204 Y2.n1203 1.1005
R11613 Y2.n86 Y2.n83 1.1005
R11614 Y2.n1169 Y2.n88 1.1005
R11615 Y2.n1170 Y2.n90 1.1005
R11616 Y2.n1172 Y2.n1171 1.1005
R11617 Y2.n1167 Y2.n1166 1.1005
R11618 Y2.n1157 Y2.n107 1.1005
R11619 Y2.n835 Y2.n834 0.733833
R11620 Y2.n703 Y2.n702 0.733833
R11621 Y2.n1334 Y2.n30 0.733833
R11622 Y2.n107 Y2.n106 0.733833
R11623 Y2.n389 Y2.n386 0.573769
R11624 Y2.n289 Y2.n286 0.573769
R11625 Y2.n759 Y2.n360 0.573695
R11626 Y2.n824 Y2.n823 0.573695
R11627 Y2.n774 Y2.n343 0.573346
R11628 Y2.n249 Y2.n247 0.550549
R11629 Y2.n1155 Y2.n110 0.550549
R11630 Y2.n394 Y2.n372 0.39244
R11631 Y2.n294 Y2.n273 0.39244
R11632 Y2.n763 Y2.n359 0.389994
R11633 Y2.n828 Y2.n261 0.389994
R11634 Y2.n779 Y2.n778 0.387191
R11635 Y2.n727 Y2.n726 0.384705
R11636 Y2.n791 Y2.n790 0.384705
R11637 Y2.n740 Y2.n388 0.384705
R11638 Y2.n804 Y2.n288 0.384705
R11639 Y2.n424 Y2.n397 0.382331
R11640 Y2.n324 Y2.n297 0.382331
R11641 Y2.n739 Y2.n395 0.382034
R11642 Y2.n803 Y2.n295 0.382034
R11643 Y2.n371 Y2.n369 0.379547
R11644 Y2.n341 Y2.n326 0.379547
R11645 Y2.n272 Y2.n269 0.379547
R11646 Y2.n764 Y2.n355 0.376968
R11647 Y2.n765 Y2.n764 0.376876
R11648 Y2.n750 Y2.n371 0.375976
R11649 Y2.n814 Y2.n272 0.375976
R11650 Y2.n339 Y2.n326 0.375884
R11651 Y2.n739 Y2.n396 0.374982
R11652 Y2.n803 Y2.n296 0.374982
R11653 Y2.n422 Y2.n397 0.374889
R11654 Y2.n322 Y2.n297 0.374889
R11655 Y2.n726 Y2.n421 0.373984
R11656 Y2.n790 Y2.n321 0.373984
R11657 Y2.n741 Y2.n740 0.373891
R11658 Y2.n805 Y2.n804 0.373891
R11659 Y2.n702 Y2.n701 0.275034
R11660 Y2.n3 Y2.n2 0.189306
R11661 Y2 Y2.n1376 0.110644
R11662 Y2.n2 Y2 0.0513955
R11663 Y2.n849 Y2.n240 0.0405
R11664 Y2.n849 Y2.n241 0.0405
R11665 Y2.n845 Y2.n241 0.0405
R11666 Y2.n845 Y2.n844 0.0405
R11667 Y2.n844 Y2.n843 0.0405
R11668 Y2.n843 Y2.n840 0.0405
R11669 Y2.n840 Y2.n198 0.0405
R11670 Y2.n942 Y2.n198 0.0405
R11671 Y2.n942 Y2.n193 0.0405
R11672 Y2.n947 Y2.n193 0.0405
R11673 Y2.n947 Y2.n196 0.0405
R11674 Y2.n196 Y2.n173 0.0405
R11675 Y2.n995 Y2.n173 0.0405
R11676 Y2.n995 Y2.n171 0.0405
R11677 Y2.n999 Y2.n154 0.0405
R11678 Y2.n1038 Y2.n154 0.0405
R11679 Y2.n1038 Y2.n151 0.0405
R11680 Y2.n1049 Y2.n151 0.0405
R11681 Y2.n1049 Y2.n152 0.0405
R11682 Y2.n1045 Y2.n152 0.0405
R11683 Y2.n1045 Y2.n1044 0.0405
R11684 Y2.n1044 Y2.n1043 0.0405
R11685 Y2.n1043 Y2.n117 0.0405
R11686 Y2.n1142 Y2.n117 0.0405
R11687 Y2.n1142 Y2.n114 0.0405
R11688 Y2.n1147 Y2.n114 0.0405
R11689 Y2.n848 Y2.n838 0.0405
R11690 Y2.n848 Y2.n847 0.0405
R11691 Y2.n847 Y2.n846 0.0405
R11692 Y2.n846 Y2.n839 0.0405
R11693 Y2.n842 Y2.n839 0.0405
R11694 Y2.n842 Y2.n841 0.0405
R11695 Y2.n841 Y2.n197 0.0405
R11696 Y2.n943 Y2.n197 0.0405
R11697 Y2.n944 Y2.n943 0.0405
R11698 Y2.n946 Y2.n944 0.0405
R11699 Y2.n946 Y2.n945 0.0405
R11700 Y2.n945 Y2.n172 0.0405
R11701 Y2.n996 Y2.n172 0.0405
R11702 Y2.n997 Y2.n996 0.0405
R11703 Y2.n998 Y2.n153 0.0405
R11704 Y2.n1039 Y2.n153 0.0405
R11705 Y2.n1040 Y2.n1039 0.0405
R11706 Y2.n1048 Y2.n1040 0.0405
R11707 Y2.n1048 Y2.n1047 0.0405
R11708 Y2.n1047 Y2.n1046 0.0405
R11709 Y2.n1046 Y2.n1041 0.0405
R11710 Y2.n1042 Y2.n1041 0.0405
R11711 Y2.n1042 Y2.n116 0.0405
R11712 Y2.n1143 Y2.n116 0.0405
R11713 Y2.n1144 Y2.n1143 0.0405
R11714 Y2.n1146 Y2.n1144 0.0405
R11715 Y2.n692 Y2.n469 0.0405
R11716 Y2.n692 Y2.n470 0.0405
R11717 Y2.n688 Y2.n470 0.0405
R11718 Y2.n688 Y2.n687 0.0405
R11719 Y2.n687 Y2.n686 0.0405
R11720 Y2.n686 Y2.n477 0.0405
R11721 Y2.n682 Y2.n477 0.0405
R11722 Y2.n682 Y2.n681 0.0405
R11723 Y2.n681 Y2.n680 0.0405
R11724 Y2.n680 Y2.n482 0.0405
R11725 Y2.n676 Y2.n482 0.0405
R11726 Y2.n676 Y2.n675 0.0405
R11727 Y2.n675 Y2.n674 0.0405
R11728 Y2.n674 Y2.n487 0.0405
R11729 Y2.n670 Y2.n669 0.0405
R11730 Y2.n669 Y2.n668 0.0405
R11731 Y2.n668 Y2.n492 0.0405
R11732 Y2.n664 Y2.n492 0.0405
R11733 Y2.n664 Y2.n663 0.0405
R11734 Y2.n663 Y2.n662 0.0405
R11735 Y2.n662 Y2.n497 0.0405
R11736 Y2.n658 Y2.n497 0.0405
R11737 Y2.n658 Y2.n657 0.0405
R11738 Y2.n657 Y2.n32 0.0405
R11739 Y2.n1344 Y2.n32 0.0405
R11740 Y2.n1344 Y2.n29 0.0405
R11741 Y2.n691 Y2.n472 0.0405
R11742 Y2.n691 Y2.n690 0.0405
R11743 Y2.n690 Y2.n689 0.0405
R11744 Y2.n689 Y2.n473 0.0405
R11745 Y2.n685 Y2.n473 0.0405
R11746 Y2.n685 Y2.n684 0.0405
R11747 Y2.n684 Y2.n683 0.0405
R11748 Y2.n683 Y2.n478 0.0405
R11749 Y2.n679 Y2.n478 0.0405
R11750 Y2.n679 Y2.n678 0.0405
R11751 Y2.n678 Y2.n677 0.0405
R11752 Y2.n677 Y2.n483 0.0405
R11753 Y2.n673 Y2.n483 0.0405
R11754 Y2.n673 Y2.n672 0.0405
R11755 Y2.n671 Y2.n488 0.0405
R11756 Y2.n667 Y2.n488 0.0405
R11757 Y2.n667 Y2.n666 0.0405
R11758 Y2.n666 Y2.n665 0.0405
R11759 Y2.n665 Y2.n493 0.0405
R11760 Y2.n661 Y2.n493 0.0405
R11761 Y2.n661 Y2.n660 0.0405
R11762 Y2.n660 Y2.n659 0.0405
R11763 Y2.n659 Y2.n498 0.0405
R11764 Y2.n498 Y2.n31 0.0405
R11765 Y2.n1345 Y2.n31 0.0405
R11766 Y2.n1346 Y2.n1345 0.0405
R11767 Y2.n999 Y2.n171 0.0360676
R11768 Y2.n998 Y2.n997 0.0360676
R11769 Y2.n670 Y2.n487 0.0360676
R11770 Y2.n672 Y2.n671 0.0360676
R11771 Y2.n276 Y2.n242 0.0360676
R11772 Y2.n279 Y2.n276 0.0360676
R11773 Y2.n280 Y2.n279 0.0360676
R11774 Y2.n281 Y2.n280 0.0360676
R11775 Y2.n282 Y2.n281 0.0360676
R11776 Y2.n303 Y2.n282 0.0360676
R11777 Y2.n314 Y2.n303 0.0360676
R11778 Y2.n315 Y2.n314 0.0360676
R11779 Y2.n316 Y2.n315 0.0360676
R11780 Y2.n317 Y2.n316 0.0360676
R11781 Y2.n333 Y2.n317 0.0360676
R11782 Y2.n334 Y2.n333 0.0360676
R11783 Y2.n335 Y2.n334 0.0360676
R11784 Y2.n349 Y2.n335 0.0360676
R11785 Y2.n350 Y2.n349 0.0360676
R11786 Y2.n351 Y2.n350 0.0360676
R11787 Y2.n375 Y2.n351 0.0360676
R11788 Y2.n376 Y2.n375 0.0360676
R11789 Y2.n379 Y2.n376 0.0360676
R11790 Y2.n380 Y2.n379 0.0360676
R11791 Y2.n381 Y2.n380 0.0360676
R11792 Y2.n382 Y2.n381 0.0360676
R11793 Y2.n403 Y2.n382 0.0360676
R11794 Y2.n414 Y2.n403 0.0360676
R11795 Y2.n415 Y2.n414 0.0360676
R11796 Y2.n416 Y2.n415 0.0360676
R11797 Y2.n417 Y2.n416 0.0360676
R11798 Y2.n433 Y2.n417 0.0360676
R11799 Y2.n434 Y2.n433 0.0360676
R11800 Y2.n435 Y2.n434 0.0360676
R11801 Y2.n452 Y2.n435 0.0360676
R11802 Y2.n453 Y2.n452 0.0360676
R11803 Y2.n454 Y2.n453 0.0360676
R11804 Y2.n277 Y2.n243 0.0360676
R11805 Y2.n278 Y2.n277 0.0360676
R11806 Y2.n278 Y2.n275 0.0360676
R11807 Y2.n810 Y2.n275 0.0360676
R11808 Y2.n810 Y2.n809 0.0360676
R11809 Y2.n809 Y2.n283 0.0360676
R11810 Y2.n313 Y2.n283 0.0360676
R11811 Y2.n313 Y2.n302 0.0360676
R11812 Y2.n796 Y2.n302 0.0360676
R11813 Y2.n796 Y2.n795 0.0360676
R11814 Y2.n795 Y2.n318 0.0360676
R11815 Y2.n784 Y2.n318 0.0360676
R11816 Y2.n784 Y2.n783 0.0360676
R11817 Y2.n783 Y2.n336 0.0360676
R11818 Y2.n770 Y2.n336 0.0360676
R11819 Y2.n770 Y2.n769 0.0360676
R11820 Y2.n769 Y2.n352 0.0360676
R11821 Y2.n377 Y2.n352 0.0360676
R11822 Y2.n378 Y2.n377 0.0360676
R11823 Y2.n378 Y2.n374 0.0360676
R11824 Y2.n746 Y2.n374 0.0360676
R11825 Y2.n746 Y2.n745 0.0360676
R11826 Y2.n745 Y2.n383 0.0360676
R11827 Y2.n413 Y2.n383 0.0360676
R11828 Y2.n413 Y2.n402 0.0360676
R11829 Y2.n732 Y2.n402 0.0360676
R11830 Y2.n732 Y2.n731 0.0360676
R11831 Y2.n731 Y2.n418 0.0360676
R11832 Y2.n720 Y2.n418 0.0360676
R11833 Y2.n720 Y2.n719 0.0360676
R11834 Y2.n719 Y2.n436 0.0360676
R11835 Y2.n706 Y2.n436 0.0360676
R11836 Y2.n706 Y2.n705 0.0360676
R11837 Y2.n1176 Y2.n95 0.0360676
R11838 Y2.n1176 Y2.n92 0.0360676
R11839 Y2.n1185 Y2.n92 0.0360676
R11840 Y2.n1185 Y2.n93 0.0360676
R11841 Y2.n1181 Y2.n93 0.0360676
R11842 Y2.n1181 Y2.n1180 0.0360676
R11843 Y2.n1180 Y2.n79 0.0360676
R11844 Y2.n1216 Y2.n79 0.0360676
R11845 Y2.n1216 Y2.n77 0.0360676
R11846 Y2.n1220 Y2.n77 0.0360676
R11847 Y2.n1220 Y2.n69 0.0360676
R11848 Y2.n1237 Y2.n69 0.0360676
R11849 Y2.n1237 Y2.n67 0.0360676
R11850 Y2.n1241 Y2.n67 0.0360676
R11851 Y2.n1241 Y2.n6 0.0360676
R11852 Y2.n1374 Y2.n6 0.0360676
R11853 Y2.n1374 Y2.n1373 0.0360676
R11854 Y2.n1373 Y2.n1372 0.0360676
R11855 Y2.n1372 Y2.n10 0.0360676
R11856 Y2.n1368 Y2.n10 0.0360676
R11857 Y2.n1368 Y2.n1367 0.0360676
R11858 Y2.n1367 Y2.n1366 0.0360676
R11859 Y2.n1366 Y2.n15 0.0360676
R11860 Y2.n1362 Y2.n15 0.0360676
R11861 Y2.n1362 Y2.n1361 0.0360676
R11862 Y2.n1361 Y2.n1360 0.0360676
R11863 Y2.n1360 Y2.n20 0.0360676
R11864 Y2.n1356 Y2.n20 0.0360676
R11865 Y2.n1356 Y2.n1355 0.0360676
R11866 Y2.n1355 Y2.n1354 0.0360676
R11867 Y2.n1354 Y2.n25 0.0360676
R11868 Y2.n1350 Y2.n25 0.0360676
R11869 Y2.n1350 Y2.n1349 0.0360676
R11870 Y2.n1177 Y2.n94 0.0360676
R11871 Y2.n1178 Y2.n1177 0.0360676
R11872 Y2.n1184 Y2.n1178 0.0360676
R11873 Y2.n1184 Y2.n1183 0.0360676
R11874 Y2.n1183 Y2.n1182 0.0360676
R11875 Y2.n1182 Y2.n1179 0.0360676
R11876 Y2.n1179 Y2.n78 0.0360676
R11877 Y2.n1217 Y2.n78 0.0360676
R11878 Y2.n1218 Y2.n1217 0.0360676
R11879 Y2.n1219 Y2.n1218 0.0360676
R11880 Y2.n1219 Y2.n68 0.0360676
R11881 Y2.n1238 Y2.n68 0.0360676
R11882 Y2.n1239 Y2.n1238 0.0360676
R11883 Y2.n1240 Y2.n1239 0.0360676
R11884 Y2.n1240 Y2.n4 0.0360676
R11885 Y2.n1375 Y2.n5 0.0360676
R11886 Y2.n1371 Y2.n5 0.0360676
R11887 Y2.n1371 Y2.n1370 0.0360676
R11888 Y2.n1370 Y2.n1369 0.0360676
R11889 Y2.n1369 Y2.n11 0.0360676
R11890 Y2.n1365 Y2.n11 0.0360676
R11891 Y2.n1365 Y2.n1364 0.0360676
R11892 Y2.n1364 Y2.n1363 0.0360676
R11893 Y2.n1363 Y2.n16 0.0360676
R11894 Y2.n1359 Y2.n16 0.0360676
R11895 Y2.n1359 Y2.n1358 0.0360676
R11896 Y2.n1358 Y2.n1357 0.0360676
R11897 Y2.n1357 Y2.n21 0.0360676
R11898 Y2.n1353 Y2.n21 0.0360676
R11899 Y2.n1353 Y2.n1352 0.0360676
R11900 Y2.n1352 Y2.n1351 0.0360676
R11901 Y2.n1351 Y2.n26 0.0360676
R11902 Y2.n1376 Y2.n1375 0.0304459
R11903 Y2.n836 Y2.n240 0.0234189
R11904 Y2.n838 Y2.n837 0.0234189
R11905 Y2.n469 Y2.n455 0.0234189
R11906 Y2.n472 Y2.n471 0.0234189
R11907 Y2.n1147 Y2.n115 0.0233108
R11908 Y2.n1146 Y2.n1145 0.0233108
R11909 Y2.n1348 Y2.n29 0.0233108
R11910 Y2.n1347 Y2.n1346 0.0233108
R11911 Y2.n837 Y2.n242 0.0227703
R11912 Y2.n836 Y2.n243 0.0227703
R11913 Y2.n115 Y2.n95 0.0227703
R11914 Y2.n1145 Y2.n94 0.0227703
R11915 Y2.n868 Y2.n867 0.0188784
R11916 Y2.n876 Y2.n875 0.0188784
R11917 Y2.n885 Y2.n884 0.0188784
R11918 Y2.n895 Y2.n894 0.0188784
R11919 Y2.n904 Y2.n903 0.0188784
R11920 Y2.n919 Y2.n199 0.0188784
R11921 Y2.n940 Y2.n201 0.0188784
R11922 Y2.n949 Y2.n192 0.0188784
R11923 Y2.n194 Y2.n189 0.0188784
R11924 Y2.n969 Y2.n182 0.0188784
R11925 Y2.n972 Y2.n971 0.0188784
R11926 Y2.n993 Y2.n175 0.0188784
R11927 Y2.n1002 Y2.n1001 0.0188784
R11928 Y2.n1015 Y2.n164 0.0188784
R11929 Y2.n1017 Y2.n155 0.0188784
R11930 Y2.n1036 Y2.n157 0.0188784
R11931 Y2.n1051 Y2.n150 0.0188784
R11932 Y2.n1065 Y2.n144 0.0188784
R11933 Y2.n1082 Y2.n1081 0.0188784
R11934 Y2.n1091 Y2.n1090 0.0188784
R11935 Y2.n1102 Y2.n1099 0.0188784
R11936 Y2.n1100 Y2.n118 0.0188784
R11937 Y2.n1140 Y2.n119 0.0188784
R11938 Y2.n542 Y2.n541 0.0188784
R11939 Y2.n546 Y2.n545 0.0188784
R11940 Y2.n550 Y2.n549 0.0188784
R11941 Y2.n554 Y2.n553 0.0188784
R11942 Y2.n559 Y2.n558 0.0188784
R11943 Y2.n571 Y2.n570 0.0188784
R11944 Y2.n576 Y2.n575 0.0188784
R11945 Y2.n583 Y2.n527 0.0188784
R11946 Y2.n586 Y2.n585 0.0188784
R11947 Y2.n590 Y2.n589 0.0188784
R11948 Y2.n595 Y2.n593 0.0188784
R11949 Y2.n603 Y2.n602 0.0188784
R11950 Y2.n607 Y2.n606 0.0188784
R11951 Y2.n611 Y2.n610 0.0188784
R11952 Y2.n615 Y2.n614 0.0188784
R11953 Y2.n622 Y2.n517 0.0188784
R11954 Y2.n625 Y2.n624 0.0188784
R11955 Y2.n630 Y2.n629 0.0188784
R11956 Y2.n643 Y2.n512 0.0188784
R11957 Y2.n646 Y2.n645 0.0188784
R11958 Y2.n648 Y2.n500 0.0188784
R11959 Y2.n655 Y2.n501 0.0188784
R11960 Y2.n507 Y2.n506 0.0188784
R11961 Y2.n835 Y2.n245 0.0188784
R11962 Y2.n266 Y2.n263 0.0188784
R11963 Y2.n821 Y2.n820 0.0188784
R11964 Y2.n817 Y2.n816 0.0188784
R11965 Y2.n767 Y2.n354 0.0188784
R11966 Y2.n365 Y2.n364 0.0188784
R11967 Y2.n757 Y2.n756 0.0188784
R11968 Y2.n753 Y2.n752 0.0188784
R11969 Y2.n1162 Y2.n106 0.0188784
R11970 Y2.n1164 Y2.n96 0.0188784
R11971 Y2.n1174 Y2.n97 0.0188784
R11972 Y2.n101 Y2.n91 0.0188784
R11973 Y2.n1257 Y2.n1256 0.0188784
R11974 Y2.n1261 Y2.n1260 0.0188784
R11975 Y2.n1268 Y2.n58 0.0188784
R11976 Y2.n1271 Y2.n1270 0.0188784
R11977 Y2.n852 Y2.n851 0.0187703
R11978 Y2.n867 Y2.n232 0.0187703
R11979 Y2.n911 Y2.n910 0.0187703
R11980 Y2.n919 Y2.n918 0.0187703
R11981 Y2.n971 Y2.n174 0.0187703
R11982 Y2.n1066 Y2.n1065 0.0187703
R11983 Y2.n1074 Y2.n1073 0.0187703
R11984 Y2.n1116 Y2.n119 0.0187703
R11985 Y2.n1118 Y2.n113 0.0187703
R11986 Y2.n694 Y2.n466 0.0187703
R11987 Y2.n541 Y2.n467 0.0187703
R11988 Y2.n562 Y2.n561 0.0187703
R11989 Y2.n570 Y2.n569 0.0187703
R11990 Y2.n595 Y2.n594 0.0187703
R11991 Y2.n631 Y2.n630 0.0187703
R11992 Y2.n634 Y2.n633 0.0187703
R11993 Y2.n506 Y2.n33 0.0187703
R11994 Y2.n1342 Y2.n34 0.0187703
R11995 Y2.n284 Y2.n274 0.0187703
R11996 Y2.n807 Y2.n285 0.0187703
R11997 Y2.n308 Y2.n306 0.0187703
R11998 Y2.n311 Y2.n309 0.0187703
R11999 Y2.n799 Y2.n798 0.0187703
R12000 Y2.n319 Y2.n301 0.0187703
R12001 Y2.n793 Y2.n320 0.0187703
R12002 Y2.n786 Y2.n331 0.0187703
R12003 Y2.n337 Y2.n332 0.0187703
R12004 Y2.n781 Y2.n338 0.0187703
R12005 Y2.n772 Y2.n346 0.0187703
R12006 Y2.n353 Y2.n348 0.0187703
R12007 Y2.n384 Y2.n373 0.0187703
R12008 Y2.n743 Y2.n385 0.0187703
R12009 Y2.n408 Y2.n406 0.0187703
R12010 Y2.n411 Y2.n409 0.0187703
R12011 Y2.n735 Y2.n734 0.0187703
R12012 Y2.n419 Y2.n401 0.0187703
R12013 Y2.n729 Y2.n420 0.0187703
R12014 Y2.n722 Y2.n431 0.0187703
R12015 Y2.n437 Y2.n432 0.0187703
R12016 Y2.n717 Y2.n438 0.0187703
R12017 Y2.n708 Y2.n449 0.0187703
R12018 Y2.n456 Y2.n451 0.0187703
R12019 Y2.n1191 Y2.n1190 0.0187703
R12020 Y2.n1195 Y2.n1194 0.0187703
R12021 Y2.n1199 Y2.n1198 0.0187703
R12022 Y2.n1201 Y2.n80 0.0187703
R12023 Y2.n1214 Y2.n81 0.0187703
R12024 Y2.n1209 Y2.n76 0.0187703
R12025 Y2.n1225 Y2.n1222 0.0187703
R12026 Y2.n1223 Y2.n70 0.0187703
R12027 Y2.n1235 Y2.n72 0.0187703
R12028 Y2.n1243 Y2.n66 0.0187703
R12029 Y2.n1250 Y2.n62 0.0187703
R12030 Y2.n1253 Y2.n1252 0.0187703
R12031 Y2.n1278 Y2.n1277 0.0187703
R12032 Y2.n1285 Y2.n54 0.0187703
R12033 Y2.n1288 Y2.n1287 0.0187703
R12034 Y2.n1293 Y2.n1292 0.0187703
R12035 Y2.n1296 Y2.n1295 0.0187703
R12036 Y2.n1305 Y2.n1304 0.0187703
R12037 Y2.n1309 Y2.n1308 0.0187703
R12038 Y2.n1313 Y2.n1312 0.0187703
R12039 Y2.n1317 Y2.n1316 0.0187703
R12040 Y2.n1324 Y2.n45 0.0187703
R12041 Y2.n1327 Y2.n1326 0.0187703
R12042 Y2.n1332 Y2.n1331 0.0187703
R12043 Y2.n875 Y2.n228 0.0185541
R12044 Y2.n1141 Y2.n118 0.0185541
R12045 Y2.n545 Y2.n538 0.0185541
R12046 Y2.n504 Y2.n501 0.0185541
R12047 Y2.n812 Y2.n811 0.0184459
R12048 Y2.n748 Y2.n747 0.0184459
R12049 Y2.n1187 Y2.n89 0.0184459
R12050 Y2.n1274 Y2.n13 0.0184459
R12051 Y2.n994 Y2.n993 0.0182297
R12052 Y2.n602 Y2.n486 0.0182297
R12053 Y2.n812 Y2.n270 0.0181216
R12054 Y2.n748 Y2.n370 0.0181216
R12055 Y2.n1187 Y2.n1186 0.0181216
R12056 Y2.n1274 Y2.n12 0.0181216
R12057 Y2.n911 Y2.n208 0.0175811
R12058 Y2.n1073 Y2.n140 0.0175811
R12059 Y2.n561 Y2.n479 0.0175811
R12060 Y2.n634 Y2.n495 0.0175811
R12061 Y2.n808 Y2.n284 0.0173649
R12062 Y2.n744 Y2.n384 0.0173649
R12063 Y2.n1191 Y2.n87 0.0173649
R12064 Y2.n1278 Y2.n14 0.0173649
R12065 Y2.n817 Y2.n268 0.0170405
R12066 Y2.n753 Y2.n368 0.0170405
R12067 Y2.n101 Y2.n100 0.0170405
R12068 Y2.n1270 Y2.n1269 0.0170405
R12069 Y2.n941 Y2.n940 0.0167162
R12070 Y2.n1051 Y2.n1050 0.0167162
R12071 Y2.n575 Y2.n480 0.0167162
R12072 Y2.n625 Y2.n494 0.0167162
R12073 Y2.n304 Y2.n285 0.0162838
R12074 Y2.n404 Y2.n385 0.0162838
R12075 Y2.n1195 Y2.n85 0.0162838
R12076 Y2.n1286 Y2.n1285 0.0162838
R12077 Y2.n970 Y2.n969 0.0159595
R12078 Y2.n1000 Y2.n164 0.0159595
R12079 Y2.n590 Y2.n485 0.0159595
R12080 Y2.n610 Y2.n489 0.0159595
R12081 Y2.n821 Y2.n267 0.0159595
R12082 Y2.n757 Y2.n367 0.0159595
R12083 Y2.n1175 Y2.n1174 0.0159595
R12084 Y2.n58 Y2.n9 0.0159595
R12085 Y2.n851 Y2.n850 0.0157432
R12086 Y2.n1118 Y2.n1117 0.0157432
R12087 Y2.n694 Y2.n693 0.0157432
R12088 Y2.n1343 Y2.n1342 0.0157432
R12089 Y2.n884 Y2.n224 0.0152027
R12090 Y2.n1102 Y2.n1101 0.0152027
R12091 Y2.n549 Y2.n474 0.0152027
R12092 Y2.n656 Y2.n500 0.0152027
R12093 Y2.n312 Y2.n308 0.0152027
R12094 Y2.n412 Y2.n408 0.0152027
R12095 Y2.n1200 Y2.n1199 0.0152027
R12096 Y2.n1288 Y2.n17 0.0152027
R12097 Y2.n1002 Y2.n170 0.0148784
R12098 Y2.n606 Y2.n522 0.0148784
R12099 Y2.n263 Y2.n262 0.0148784
R12100 Y2.n364 Y2.n363 0.0148784
R12101 Y2.n1164 Y2.n1163 0.0148784
R12102 Y2.n1260 Y2.n8 0.0148784
R12103 Y2.n904 Y2.n212 0.0141216
R12104 Y2.n1081 Y2.n135 0.0141216
R12105 Y2.n560 Y2.n559 0.0141216
R12106 Y2.n512 Y2.n496 0.0141216
R12107 Y2.n309 Y2.n300 0.0141216
R12108 Y2.n409 Y2.n400 0.0141216
R12109 Y2.n1215 Y2.n80 0.0141216
R12110 Y2.n1293 Y2.n18 0.0141216
R12111 Y2.n471 Y2.n454 0.0137973
R12112 Y2.n705 Y2.n455 0.0137973
R12113 Y2.n768 Y2.n767 0.0137973
R12114 Y2.n704 Y2.n703 0.0137973
R12115 Y2.n1256 Y2.n7 0.0137973
R12116 Y2.n30 Y2.n28 0.0137973
R12117 Y2.n1349 Y2.n1348 0.0137973
R12118 Y2.n1347 Y2.n26 0.0137973
R12119 Y2.n1335 Y2.n40 0.0134381
R12120 Y2.n200 Y2.n192 0.0133649
R12121 Y2.n157 Y2.n156 0.0133649
R12122 Y2.n527 Y2.n481 0.0133649
R12123 Y2.n623 Y2.n622 0.0133649
R12124 Y2.n798 Y2.n797 0.0130405
R12125 Y2.n734 Y2.n733 0.0130405
R12126 Y2.n1208 Y2.n81 0.0130405
R12127 Y2.n1295 Y2.n19 0.0130405
R12128 Y2.n771 Y2.n348 0.0128243
R12129 Y2.n707 Y2.n451 0.0128243
R12130 Y2.n1252 Y2.n1251 0.0128243
R12131 Y2.n1331 Y2.n27 0.0128243
R12132 Y2.n195 Y2.n194 0.0126081
R12133 Y2.n1017 Y2.n1016 0.0126081
R12134 Y2.n586 Y2.n484 0.0126081
R12135 Y2.n614 Y2.n490 0.0126081
R12136 Y2.n244 Y2.n239 0.0123919
R12137 Y2.n1149 Y2.n1148 0.0123919
R12138 Y2.n468 Y2.n457 0.0123919
R12139 Y2.n42 Y2.n41 0.0123919
R12140 Y2.n794 Y2.n319 0.0119595
R12141 Y2.n730 Y2.n419 0.0119595
R12142 Y2.n1221 Y2.n76 0.0119595
R12143 Y2.n1305 Y2.n50 0.0119595
R12144 Y2.n894 Y2.n220 0.0118514
R12145 Y2.n1091 Y2.n126 0.0118514
R12146 Y2.n553 Y2.n475 0.0118514
R12147 Y2.n646 Y2.n499 0.0118514
R12148 Y2.n346 Y2.n345 0.0117432
R12149 Y2.n449 Y2.n448 0.0117432
R12150 Y2.n1242 Y2.n62 0.0117432
R12151 Y2.n1326 Y2.n1325 0.0117432
R12152 Y2.n701 Y2.n698 0.0116588
R12153 Y2.n835 Y2.n244 0.011527
R12154 Y2.n703 Y2.n457 0.011527
R12155 Y2.n1149 Y2.n106 0.0114189
R12156 Y2.n42 Y2.n30 0.0114189
R12157 Y2.n1171 Y2.n1170 0.0109762
R12158 Y2.n1169 Y2.n83 0.0109762
R12159 Y2.n1205 Y2.n1204 0.0109762
R12160 Y2.n1228 Y2.n74 0.0109762
R12161 Y2.n1229 Y2.n64 0.0109762
R12162 Y2.n1247 Y2.n1246 0.0109762
R12163 Y2.n1264 Y2.n60 0.0109762
R12164 Y2.n1265 Y2.n56 0.0109762
R12165 Y2.n1282 Y2.n1281 0.0109762
R12166 Y2.n1299 Y2.n52 0.0109762
R12167 Y2.n1301 Y2.n1300 0.0109762
R12168 Y2.n1320 Y2.n47 0.0109762
R12169 Y2.n1321 Y2.n40 0.0109762
R12170 Y2.n697 Y2.n462 0.0109762
R12171 Y2.n536 Y2.n462 0.0109762
R12172 Y2.n536 Y2.n535 0.0109762
R12173 Y2.n535 Y2.n532 0.0109762
R12174 Y2.n565 Y2.n532 0.0109762
R12175 Y2.n566 Y2.n565 0.0109762
R12176 Y2.n566 Y2.n529 0.0109762
R12177 Y2.n579 Y2.n529 0.0109762
R12178 Y2.n580 Y2.n579 0.0109762
R12179 Y2.n580 Y2.n524 0.0109762
R12180 Y2.n598 Y2.n524 0.0109762
R12181 Y2.n600 Y2.n599 0.0109762
R12182 Y2.n599 Y2.n519 0.0109762
R12183 Y2.n618 Y2.n519 0.0109762
R12184 Y2.n619 Y2.n618 0.0109762
R12185 Y2.n619 Y2.n514 0.0109762
R12186 Y2.n637 Y2.n514 0.0109762
R12187 Y2.n638 Y2.n637 0.0109762
R12188 Y2.n638 Y2.n510 0.0109762
R12189 Y2.n651 Y2.n510 0.0109762
R12190 Y2.n652 Y2.n651 0.0109762
R12191 Y2.n652 Y2.n37 0.0109762
R12192 Y2.n1339 Y2.n37 0.0109762
R12193 Y2.n272 Y2.n271 0.0109762
R12194 Y2.n804 Y2.n294 0.0109762
R12195 Y2.n803 Y2.n802 0.0109762
R12196 Y2.n790 Y2.n297 0.0109762
R12197 Y2.n789 Y2.n326 0.0109762
R12198 Y2.n778 Y2.n344 0.0109762
R12199 Y2.n764 Y2.n763 0.0109762
R12200 Y2.n371 Y2.n361 0.0109762
R12201 Y2.n740 Y2.n394 0.0109762
R12202 Y2.n739 Y2.n738 0.0109762
R12203 Y2.n726 Y2.n397 0.0109762
R12204 Y2.n1170 Y2.n1169 0.01095
R12205 Y2.n1204 Y2.n83 0.01095
R12206 Y2.n1205 Y2.n74 0.01095
R12207 Y2.n1229 Y2.n1228 0.01095
R12208 Y2.n1246 Y2.n64 0.01095
R12209 Y2.n1247 Y2.n60 0.01095
R12210 Y2.n1265 Y2.n1264 0.01095
R12211 Y2.n1281 Y2.n56 0.01095
R12212 Y2.n1282 Y2.n52 0.01095
R12213 Y2.n1301 Y2.n1299 0.01095
R12214 Y2.n1300 Y2.n47 0.01095
R12215 Y2.n1321 Y2.n1320 0.01095
R12216 Y2.n600 Y2.n598 0.01095
R12217 Y2.n1339 Y2.n1338 0.01095
R12218 Y2.n271 Y2.n261 0.01095
R12219 Y2.n294 Y2.n272 0.01095
R12220 Y2.n804 Y2.n803 0.01095
R12221 Y2.n802 Y2.n297 0.01095
R12222 Y2.n790 Y2.n789 0.01095
R12223 Y2.n778 Y2.n326 0.01095
R12224 Y2.n764 Y2.n344 0.01095
R12225 Y2.n763 Y2.n361 0.01095
R12226 Y2.n394 Y2.n371 0.01095
R12227 Y2.n740 Y2.n739 0.01095
R12228 Y2.n738 Y2.n397 0.01095
R12229 Y2.n726 Y2.n725 0.01095
R12230 Y2.n330 Y2.n320 0.0108784
R12231 Y2.n430 Y2.n420 0.0108784
R12232 Y2.n1225 Y2.n1224 0.0108784
R12233 Y2.n1309 Y2.n22 0.0108784
R12234 Y2.n895 Y2.n216 0.0107703
R12235 Y2.n1090 Y2.n130 0.0107703
R12236 Y2.n554 Y2.n476 0.0107703
R12237 Y2.n645 Y2.n644 0.0107703
R12238 Y2.n782 Y2.n781 0.0106622
R12239 Y2.n718 Y2.n717 0.0106622
R12240 Y2.n71 Y2.n66 0.0106622
R12241 Y2.n45 Y2.n24 0.0106622
R12242 Y2.n698 Y2.n697 0.0106095
R12243 Y2.n948 Y2.n189 0.0100135
R12244 Y2.n1037 Y2.n155 0.0100135
R12245 Y2.n585 Y2.n584 0.0100135
R12246 Y2.n615 Y2.n491 0.0100135
R12247 Y2.n786 Y2.n785 0.0097973
R12248 Y2.n722 Y2.n721 0.0097973
R12249 Y2.n1236 Y2.n70 0.0097973
R12250 Y2.n1313 Y2.n23 0.0097973
R12251 Y2.n701 Y2.n700 0.00967266
R12252 Y2.n785 Y2.n332 0.00958108
R12253 Y2.n721 Y2.n432 0.00958108
R12254 Y2.n1236 Y2.n1235 0.00958108
R12255 Y2.n1316 Y2.n23 0.00958108
R12256 Y2.n949 Y2.n948 0.00925676
R12257 Y2.n1037 Y2.n1036 0.00925676
R12258 Y2.n584 Y2.n583 0.00925676
R12259 Y2.n517 Y2.n491 0.00925676
R12260 Y2.n778 Y2.n343 0.00880612
R12261 Y2.n782 Y2.n337 0.00871622
R12262 Y2.n718 Y2.n437 0.00871622
R12263 Y2.n72 Y2.n71 0.00871622
R12264 Y2.n1317 Y2.n24 0.00871622
R12265 Y2.n903 Y2.n216 0.0085
R12266 Y2.n1082 Y2.n130 0.0085
R12267 Y2.n558 Y2.n476 0.0085
R12268 Y2.n644 Y2.n643 0.0085
R12269 Y2.n331 Y2.n330 0.0085
R12270 Y2.n431 Y2.n430 0.0085
R12271 Y2.n1224 Y2.n1223 0.0085
R12272 Y2.n1312 Y2.n22 0.0085
R12273 Y2.n1171 Y2.n1168 0.00809524
R12274 Y2.n699 Y2.n447 0.00778095
R12275 Y2.n345 Y2.n338 0.00763514
R12276 Y2.n448 Y2.n438 0.00763514
R12277 Y2.n1243 Y2.n1242 0.00763514
R12278 Y2.n1325 Y2.n1324 0.00763514
R12279 Y2.n885 Y2.n220 0.00741892
R12280 Y2.n1099 Y2.n126 0.00741892
R12281 Y2.n550 Y2.n475 0.00741892
R12282 Y2.n648 Y2.n499 0.00741892
R12283 Y2.n794 Y2.n793 0.00741892
R12284 Y2.n730 Y2.n729 0.00741892
R12285 Y2.n1222 Y2.n1221 0.00741892
R12286 Y2.n1308 Y2.n50 0.00741892
R12287 Y2.n725 Y2.n426 0.00725714
R12288 Y2.n700 Y2.n699 0.00707381
R12289 Y2.n852 Y2.n239 0.00698649
R12290 Y2.n1148 Y2.n113 0.00698649
R12291 Y2.n468 Y2.n466 0.00698649
R12292 Y2.n41 Y2.n34 0.00698649
R12293 Y2.n831 Y2.n261 0.00696162
R12294 Y2.n1338 Y2.n38 0.00691667
R12295 Y2.n195 Y2.n182 0.00666216
R12296 Y2.n1016 Y2.n1015 0.00666216
R12297 Y2.n589 Y2.n484 0.00666216
R12298 Y2.n611 Y2.n490 0.00666216
R12299 Y2.n772 Y2.n771 0.00655405
R12300 Y2.n708 Y2.n707 0.00655405
R12301 Y2.n1251 Y2.n1250 0.00655405
R12302 Y2.n1327 Y2.n27 0.00655405
R12303 Y2.n797 Y2.n301 0.00633784
R12304 Y2.n733 Y2.n401 0.00633784
R12305 Y2.n1209 Y2.n1208 0.00633784
R12306 Y2.n1304 Y2.n19 0.00633784
R12307 Y2.n1376 Y2.n4 0.00612162
R12308 Y2.n201 Y2.n200 0.00590541
R12309 Y2.n156 Y2.n150 0.00590541
R12310 Y2.n576 Y2.n481 0.00590541
R12311 Y2.n624 Y2.n623 0.00590541
R12312 Y2.n763 Y2.n360 0.00588776
R12313 Y2.n824 Y2.n261 0.00588776
R12314 Y2.n768 Y2.n353 0.00547297
R12315 Y2.n704 Y2.n456 0.00547297
R12316 Y2.n1253 Y2.n7 0.00547297
R12317 Y2.n1332 Y2.n28 0.00547297
R12318 Y2.n799 Y2.n300 0.00525676
R12319 Y2.n735 Y2.n400 0.00525676
R12320 Y2.n1215 Y2.n1214 0.00525676
R12321 Y2.n1296 Y2.n18 0.00525676
R12322 Y2.n910 Y2.n212 0.00514865
R12323 Y2.n1074 Y2.n135 0.00514865
R12324 Y2.n562 Y2.n560 0.00514865
R12325 Y2.n633 Y2.n496 0.00514865
R12326 Y2.n1336 Y2.n1335 0.00440238
R12327 Y2.n175 Y2.n170 0.00439189
R12328 Y2.n603 Y2.n522 0.00439189
R12329 Y2.n262 Y2.n245 0.00439189
R12330 Y2.n363 Y2.n354 0.00439189
R12331 Y2.n1163 Y2.n1162 0.00439189
R12332 Y2.n1257 Y2.n8 0.00439189
R12333 Y2.n464 Y2.n463 0.00425921
R12334 Y2.n695 Y2.n465 0.00425921
R12335 Y2.n555 Y2.n552 0.00425921
R12336 Y2.n557 Y2.n533 0.00425921
R12337 Y2.n572 Y2.n530 0.00425921
R12338 Y2.n577 Y2.n574 0.00425921
R12339 Y2.n582 Y2.n528 0.00425921
R12340 Y2.n587 Y2.n526 0.00425921
R12341 Y2.n604 Y2.n601 0.00425921
R12342 Y2.n616 Y2.n613 0.00425921
R12343 Y2.n621 Y2.n518 0.00425921
R12344 Y2.n626 Y2.n516 0.00425921
R12345 Y2.n628 Y2.n515 0.00425921
R12346 Y2.n642 Y2.n640 0.00425921
R12347 Y2.n647 Y2.n511 0.00425921
R12348 Y2.n1341 Y2.n35 0.00425921
R12349 Y2.n43 Y2.n36 0.00425921
R12350 Y2.n328 Y2.n327 0.00425921
R12351 Y2.n787 Y2.n329 0.00425921
R12352 Y2.n428 Y2.n427 0.00425921
R12353 Y2.n723 Y2.n429 0.00425921
R12354 Y2.n102 Y2.n99 0.00425921
R12355 Y2.n1189 Y2.n1188 0.00425921
R12356 Y2.n1193 Y2.n1192 0.00425921
R12357 Y2.n1197 Y2.n1196 0.00425921
R12358 Y2.n1207 Y2.n75 0.00425921
R12359 Y2.n1226 Y2.n73 0.00425921
R12360 Y2.n1234 Y2.n1231 0.00425921
R12361 Y2.n1232 Y2.n65 0.00425921
R12362 Y2.n1258 Y2.n1255 0.00425921
R12363 Y2.n1272 Y2.n57 0.00425921
R12364 Y2.n1276 Y2.n1275 0.00425921
R12365 Y2.n1279 Y2.n55 0.00425921
R12366 Y2.n1284 Y2.n53 0.00425921
R12367 Y2.n1307 Y2.n1306 0.00425921
R12368 Y2.n1311 Y2.n1310 0.00425921
R12369 Y2.n1315 Y2.n1314 0.00425921
R12370 Y2.n1318 Y2.n46 0.00425921
R12371 Y2.n446 Y2.n445 0.00424524
R12372 Y2.n540 Y2.n465 0.0042371
R12373 Y2.n544 Y2.n543 0.0042371
R12374 Y2.n548 Y2.n547 0.0042371
R12375 Y2.n552 Y2.n551 0.0042371
R12376 Y2.n563 Y2.n531 0.0042371
R12377 Y2.n568 Y2.n530 0.0042371
R12378 Y2.n588 Y2.n587 0.0042371
R12379 Y2.n592 Y2.n591 0.0042371
R12380 Y2.n596 Y2.n523 0.0042371
R12381 Y2.n601 Y2.n523 0.0042371
R12382 Y2.n605 Y2.n604 0.0042371
R12383 Y2.n609 Y2.n608 0.0042371
R12384 Y2.n613 Y2.n612 0.0042371
R12385 Y2.n632 Y2.n515 0.0042371
R12386 Y2.n635 Y2.n513 0.0042371
R12387 Y2.n649 Y2.n647 0.0042371
R12388 Y2.n654 Y2.n502 0.0042371
R12389 Y2.n509 Y2.n508 0.0042371
R12390 Y2.n505 Y2.n35 0.0042371
R12391 Y2.n819 Y2.n818 0.0042371
R12392 Y2.n310 Y2.n298 0.0042371
R12393 Y2.n800 Y2.n299 0.0042371
R12394 Y2.n357 Y2.n356 0.0042371
R12395 Y2.n755 Y2.n754 0.0042371
R12396 Y2.n410 Y2.n398 0.0042371
R12397 Y2.n736 Y2.n399 0.0042371
R12398 Y2.n710 Y2.n709 0.0042371
R12399 Y2.n460 Y2.n459 0.0042371
R12400 Y2.n1173 Y2.n98 0.0042371
R12401 Y2.n103 Y2.n102 0.0042371
R12402 Y2.n1197 Y2.n84 0.0042371
R12403 Y2.n1202 Y2.n82 0.0042371
R12404 Y2.n1213 Y2.n1212 0.0042371
R12405 Y2.n1210 Y2.n1207 0.0042371
R12406 Y2.n1244 Y2.n65 0.0042371
R12407 Y2.n1249 Y2.n63 0.0042371
R12408 Y2.n1254 Y2.n61 0.0042371
R12409 Y2.n1255 Y2.n1254 0.0042371
R12410 Y2.n1259 Y2.n1258 0.0042371
R12411 Y2.n1262 Y2.n59 0.0042371
R12412 Y2.n1267 Y2.n57 0.0042371
R12413 Y2.n1289 Y2.n53 0.0042371
R12414 Y2.n1294 Y2.n1291 0.0042371
R12415 Y2.n1297 Y2.n51 0.0042371
R12416 Y2.n1306 Y2.n1303 0.0042371
R12417 Y2.n1323 Y2.n46 0.0042371
R12418 Y2.n1328 Y2.n44 0.0042371
R12419 Y2.n1333 Y2.n1330 0.0042371
R12420 Y2.n1334 Y2.n1333 0.0042371
R12421 Y2.n1159 Y2.n1157 0.00423273
R12422 Y2.n260 Y2.n259 0.00422178
R12423 Y2.n1156 Y2.n108 0.00422178
R12424 Y2.n444 Y2.n426 0.00421905
R12425 Y2.n312 Y2.n311 0.00417568
R12426 Y2.n412 Y2.n411 0.00417568
R12427 Y2.n1201 Y2.n1200 0.00417568
R12428 Y2.n1292 Y2.n17 0.00417568
R12429 Y2.n543 Y2.n539 0.00410442
R12430 Y2.n508 Y2.n503 0.00410442
R12431 Y2.n876 Y2.n224 0.00406757
R12432 Y2.n1101 Y2.n1100 0.00406757
R12433 Y2.n546 Y2.n474 0.00406757
R12434 Y2.n656 Y2.n655 0.00406757
R12435 Y2.n774 Y2.n773 0.00402269
R12436 Y2.n813 Y2.n273 0.00398793
R12437 Y2.n749 Y2.n372 0.00398793
R12438 Y2.n1188 Y2.n90 0.00397174
R12439 Y2.n1234 Y2.n1233 0.00397174
R12440 Y2.n1275 Y2.n1273 0.00397174
R12441 Y2.n1319 Y2.n1315 0.00397174
R12442 Y2.n582 Y2.n581 0.00394963
R12443 Y2.n617 Y2.n518 0.00394963
R12444 Y2.n823 Y2.n822 0.00394626
R12445 Y2.n759 Y2.n758 0.00394626
R12446 Y2.n829 Y2.n828 0.00393696
R12447 Y2.n359 Y2.n358 0.00393696
R12448 Y2.n806 Y2.n286 0.00390294
R12449 Y2.n742 Y2.n386 0.00390294
R12450 Y2.n780 Y2.n779 0.00389381
R12451 Y2.n305 Y2.n288 0.00385851
R12452 Y2.n791 Y2.n325 0.00385851
R12453 Y2.n405 Y2.n388 0.00385851
R12454 Y2.n727 Y2.n425 0.00385851
R12455 Y2.n305 Y2.n295 0.00380768
R12456 Y2.n405 Y2.n395 0.00380768
R12457 Y2.n325 Y2.n324 0.00380053
R12458 Y2.n425 Y2.n424 0.00380053
R12459 Y2.n557 Y2.n556 0.00379484
R12460 Y2.n642 Y2.n641 0.00379484
R12461 Y2.n1160 Y2.n107 0.00379484
R12462 Y2.n702 Y2.n461 0.00377273
R12463 Y2.n818 Y2.n269 0.0037725
R12464 Y2.n780 Y2.n341 0.0037725
R12465 Y2.n754 Y2.n369 0.0037725
R12466 Y2.n714 Y2.n713 0.00374762
R12467 Y2.n358 Y2.n355 0.00372958
R12468 Y2.n1203 Y2.n1202 0.0037285
R12469 Y2.n1291 Y2.n1290 0.0037285
R12470 Y2.n765 Y2.n357 0.00372177
R12471 Y2.n1212 Y2.n1211 0.00370639
R12472 Y2.n1302 Y2.n51 0.00370639
R12473 Y2.n712 Y2.n447 0.00369524
R12474 Y2.n567 Y2.n531 0.00366216
R12475 Y2.n636 Y2.n635 0.00366216
R12476 Y2.n441 Y2.n439 0.00366216
R12477 Y2.n443 Y2.n442 0.00364005
R12478 Y2.n850 Y2.n232 0.00363514
R12479 Y2.n1117 Y2.n1116 0.00363514
R12480 Y2.n693 Y2.n467 0.00363514
R12481 Y2.n1343 Y2.n33 0.00363514
R12482 Y2.n1158 Y2.n104 0.00359048
R12483 Y2.n339 Y2.n329 0.00358532
R12484 Y2.n259 Y2.n249 0.00357902
R12485 Y2.n110 Y2.n108 0.00357902
R12486 Y2.n814 Y2.n813 0.00357098
R12487 Y2.n750 Y2.n749 0.00357098
R12488 Y2.n574 Y2.n573 0.00348526
R12489 Y2.n627 Y2.n626 0.00348526
R12490 Y2.n310 Y2.n296 0.003457
R12491 Y2.n410 Y2.n396 0.003457
R12492 Y2.n322 Y2.n299 0.00344926
R12493 Y2.n422 Y2.n399 0.00344926
R12494 Y2.n1193 Y2.n86 0.00344103
R12495 Y2.n1227 Y2.n1226 0.00344103
R12496 Y2.n1283 Y2.n55 0.00344103
R12497 Y2.n1310 Y2.n49 0.00344103
R12498 Y2.n792 Y2.n321 0.00343273
R12499 Y2.n728 Y2.n421 0.00343273
R12500 Y2.n805 Y2.n287 0.00341839
R12501 Y2.n741 Y2.n387 0.00341839
R12502 Y2.n394 Y2.n389 0.00341837
R12503 Y2.n294 Y2.n289 0.00341837
R12504 Y2.n1168 Y2.n1167 0.00335476
R12505 Y2.n548 Y2.n534 0.00335258
R12506 Y2.n650 Y2.n502 0.00335258
R12507 Y2.n806 Y2.n805 0.0033136
R12508 Y2.n742 Y2.n741 0.0033136
R12509 Y2.n972 Y2.n970 0.00331081
R12510 Y2.n1001 Y2.n1000 0.00331081
R12511 Y2.n593 Y2.n485 0.00331081
R12512 Y2.n607 Y2.n489 0.00331081
R12513 Y2.n267 Y2.n266 0.00331081
R12514 Y2.n367 Y2.n365 0.00331081
R12515 Y2.n1175 Y2.n96 0.00331081
R12516 Y2.n1261 Y2.n9 0.00331081
R12517 Y2.n323 Y2.n322 0.00330444
R12518 Y2.n423 Y2.n422 0.00330444
R12519 Y2.n327 Y2.n321 0.0032992
R12520 Y2.n427 Y2.n421 0.0032992
R12521 Y2.n307 Y2.n296 0.00329663
R12522 Y2.n407 Y2.n396 0.00329663
R12523 Y2.n715 Y2.n440 0.00324201
R12524 Y2.n591 Y2.n525 0.00319779
R12525 Y2.n609 Y2.n520 0.00319779
R12526 Y2.n711 Y2.n710 0.00319779
R12527 Y2.n1245 Y2.n63 0.00319779
R12528 Y2.n1322 Y2.n44 0.00319779
R12529 Y2.n822 Y2.n265 0.00317568
R12530 Y2.n758 Y2.n366 0.00317568
R12531 Y2.n1173 Y2.n1172 0.00317568
R12532 Y2.n1266 Y2.n59 0.00317568
R12533 Y2.n815 Y2.n814 0.00316007
R12534 Y2.n751 Y2.n750 0.00316007
R12535 Y2.n340 Y2.n339 0.00314581
R12536 Y2.n1165 Y2.n105 0.00310934
R12537 Y2.n306 Y2.n304 0.00309459
R12538 Y2.n406 Y2.n404 0.00309459
R12539 Y2.n1198 Y2.n85 0.00309459
R12540 Y2.n1287 Y2.n1286 0.00309459
R12541 Y2.n696 Y2.n464 0.003043
R12542 Y2.n1340 Y2.n36 0.003043
R12543 Y2.n766 Y2.n355 0.00302306
R12544 Y2.n766 Y2.n765 0.00300884
R12545 Y2.n881 Y2.n879 0.0029881
R12546 Y2.n914 Y2.n210 0.0029881
R12547 Y2.n937 Y2.n929 0.0029881
R12548 Y2.n1055 Y2.n1054 0.0029881
R12549 Y2.n341 Y2.n340 0.00298054
R12550 Y2.n815 Y2.n269 0.00298054
R12551 Y2.n751 Y2.n369 0.00298054
R12552 Y2.n1070 Y2.n138 0.0029619
R12553 Y2.n1105 Y2.n124 0.0029619
R12554 Y2.n324 Y2.n323 0.00293083
R12555 Y2.n424 Y2.n423 0.00293083
R12556 Y2.n307 Y2.n295 0.0029237
R12557 Y2.n407 Y2.n395 0.0029237
R12558 Y2.n597 Y2.n592 0.00291032
R12559 Y2.n608 Y2.n521 0.00291032
R12560 Y2.n773 Y2.n347 0.00291032
R12561 Y2.n709 Y2.n450 0.00291032
R12562 Y2.n1166 Y2.n98 0.00291032
R12563 Y2.n1249 Y2.n1248 0.00291032
R12564 Y2.n1263 Y2.n1262 0.00291032
R12565 Y2.n1329 Y2.n1328 0.00291032
R12566 Y2.n288 Y2.n287 0.00289527
R12567 Y2.n388 Y2.n387 0.00289527
R12568 Y2.n792 Y2.n791 0.00289527
R12569 Y2.n728 Y2.n727 0.00289527
R12570 Y2.n257 Y2.n249 0.00287188
R12571 Y2.n1153 Y2.n110 0.00284569
R12572 Y2.n779 Y2.n342 0.00283826
R12573 Y2.n1336 Y2.n38 0.00283095
R12574 Y2.n828 Y2.n827 0.00279542
R12575 Y2.n362 Y2.n359 0.00279542
R12576 Y2.n290 Y2.n273 0.00276679
R12577 Y2.n390 Y2.n372 0.00276679
R12578 Y2.n547 Y2.n537 0.00275553
R12579 Y2.n654 Y2.n653 0.00275553
R12580 Y2.n463 Y2.n458 0.00273342
R12581 Y2.n1334 Y2.n43 0.00273342
R12582 Y2.n257 Y2.n256 0.00272619
R12583 Y2.n256 Y2.n255 0.00272619
R12584 Y2.n855 Y2.n237 0.00272619
R12585 Y2.n857 Y2.n856 0.00272619
R12586 Y2.n865 Y2.n864 0.00272619
R12587 Y2.n873 Y2.n226 0.00272619
R12588 Y2.n878 Y2.n226 0.00272619
R12589 Y2.n880 Y2.n222 0.00272619
R12590 Y2.n888 Y2.n222 0.00272619
R12591 Y2.n890 Y2.n218 0.00272619
R12592 Y2.n898 Y2.n218 0.00272619
R12593 Y2.n906 Y2.n214 0.00272619
R12594 Y2.n907 Y2.n906 0.00272619
R12595 Y2.n916 Y2.n915 0.00272619
R12596 Y2.n916 Y2.n206 0.00272619
R12597 Y2.n924 Y2.n204 0.00272619
R12598 Y2.n928 Y2.n204 0.00272619
R12599 Y2.n936 Y2.n935 0.00272619
R12600 Y2.n931 Y2.n930 0.00272619
R12601 Y2.n954 Y2.n187 0.00272619
R12602 Y2.n964 Y2.n963 0.00272619
R12603 Y2.n967 Y2.n964 0.00272619
R12604 Y2.n975 Y2.n180 0.00272619
R12605 Y2.n976 Y2.n975 0.00272619
R12606 Y2.n977 Y2.n976 0.00272619
R12607 Y2.n991 Y2.n990 0.00272619
R12608 Y2.n1005 Y2.n168 0.00272619
R12609 Y2.n1006 Y2.n1005 0.00272619
R12610 Y2.n1012 Y2.n1011 0.00272619
R12611 Y2.n1013 Y2.n1012 0.00272619
R12612 Y2.n1013 Y2.n162 0.00272619
R12613 Y2.n1022 Y2.n160 0.00272619
R12614 Y2.n1026 Y2.n160 0.00272619
R12615 Y2.n1032 Y2.n1031 0.00272619
R12616 Y2.n1031 Y2.n1028 0.00272619
R12617 Y2.n1060 Y2.n146 0.00272619
R12618 Y2.n1069 Y2.n1068 0.00272619
R12619 Y2.n1077 Y2.n1076 0.00272619
R12620 Y2.n1079 Y2.n1078 0.00272619
R12621 Y2.n1088 Y2.n1087 0.00272619
R12622 Y2.n1097 Y2.n1096 0.00272619
R12623 Y2.n1096 Y2.n124 0.00272619
R12624 Y2.n1107 Y2.n1106 0.00272619
R12625 Y2.n1107 Y2.n122 0.00272619
R12626 Y2.n1111 Y2.n122 0.00272619
R12627 Y2.n1136 Y2.n1135 0.00272619
R12628 Y2.n1135 Y2.n1113 0.00272619
R12629 Y2.n1126 Y2.n1115 0.00272619
R12630 Y2.n1126 Y2.n1125 0.00272619
R12631 Y2.n1152 Y2.n111 0.00272619
R12632 Y2.n1154 Y2.n1153 0.00272619
R12633 Y2.n255 Y2.n254 0.0027
R12634 Y2.n856 Y2.n855 0.0027
R12635 Y2.n865 Y2.n863 0.0027
R12636 Y2.n873 Y2.n872 0.0027
R12637 Y2.n881 Y2.n880 0.0027
R12638 Y2.n908 Y2.n907 0.0027
R12639 Y2.n935 Y2.n930 0.0027
R12640 Y2.n954 Y2.n953 0.0027
R12641 Y2.n963 Y2.n185 0.0027
R12642 Y2.n991 Y2.n983 0.0027
R12643 Y2.n984 Y2.n168 0.0027
R12644 Y2.n1028 Y2.n148 0.0027
R12645 Y2.n1056 Y2.n146 0.0027
R12646 Y2.n1068 Y2.n142 0.0027
R12647 Y2.n1079 Y2.n1077 0.0027
R12648 Y2.n1088 Y2.n1086 0.0027
R12649 Y2.n1097 Y2.n1095 0.0027
R12650 Y2.n1125 Y2.n1124 0.0027
R12651 Y2.n1154 Y2.n1152 0.0027
R12652 Y2.n908 Y2.n210 0.00264762
R12653 Y2.n1076 Y2.n138 0.00264762
R12654 Y2.n1192 Y2.n88 0.00264496
R12655 Y2.n1280 Y2.n1279 0.00264496
R12656 Y2.n788 Y2.n328 0.00262285
R12657 Y2.n724 Y2.n428 0.00262285
R12658 Y2.n1230 Y2.n73 0.00262285
R12659 Y2.n1311 Y2.n48 0.00262285
R12660 Y2.n929 Y2.n928 0.00262143
R12661 Y2.n1056 Y2.n1055 0.00262143
R12662 Y2.n578 Y2.n577 0.00260074
R12663 Y2.n620 Y2.n516 0.00260074
R12664 Y2.n883 Y2.n225 0.00257862
R12665 Y2.n1104 Y2.n1103 0.00257862
R12666 Y2.n1054 Y2.n148 0.00256905
R12667 Y2.n941 Y2.n199 0.00255405
R12668 Y2.n1050 Y2.n144 0.00255405
R12669 Y2.n571 Y2.n480 0.00255405
R12670 Y2.n629 Y2.n494 0.00255405
R12671 Y2.n937 Y2.n936 0.00254286
R12672 Y2.n1070 Y2.n1069 0.00254286
R12673 Y2.n939 Y2.n938 0.0025344
R12674 Y2.n915 Y2.n914 0.00251667
R12675 Y2.n1053 Y2.n1052 0.00251228
R12676 Y2.n833 Y2.n832 0.0024936
R12677 Y2.n879 Y2.n878 0.00246429
R12678 Y2.n1106 Y2.n1105 0.00246429
R12679 Y2.n564 Y2.n563 0.00244595
R12680 Y2.n639 Y2.n513 0.00244595
R12681 Y2.n899 Y2.n898 0.0024381
R12682 Y2.n1086 Y2.n1085 0.0024381
R12683 Y2.n912 Y2.n211 0.00242383
R12684 Y2.n1072 Y2.n139 0.00242383
R12685 Y2.n1159 Y2.n1158 0.00238571
R12686 Y2.n714 Y2.n446 0.00238571
R12687 Y2.n862 Y2.n235 0.00238571
R12688 Y2.n871 Y2.n230 0.00238571
R12689 Y2.n891 Y2.n889 0.00238571
R12690 Y2.n900 Y2.n899 0.00238571
R12691 Y2.n923 Y2.n922 0.00238571
R12692 Y2.n952 Y2.n190 0.00238571
R12693 Y2.n959 Y2.n958 0.00238571
R12694 Y2.n982 Y2.n178 0.00238571
R12695 Y2.n989 Y2.n985 0.00238571
R12696 Y2.n1007 Y2.n1006 0.00238571
R12697 Y2.n1021 Y2.n1020 0.00238571
R12698 Y2.n1033 Y2.n1027 0.00238571
R12699 Y2.n1062 Y2.n1061 0.00238571
R12700 Y2.n1085 Y2.n133 0.00238571
R12701 Y2.n1094 Y2.n128 0.00238571
R12702 Y2.n1137 Y2.n1112 0.00238571
R12703 Y2.n1131 Y2.n1130 0.00238571
R12704 Y2.n854 Y2.n853 0.00237961
R12705 Y2.n858 Y2.n236 0.00237961
R12706 Y2.n866 Y2.n234 0.00237961
R12707 Y2.n874 Y2.n227 0.00237961
R12708 Y2.n877 Y2.n227 0.00237961
R12709 Y2.n886 Y2.n223 0.00237961
R12710 Y2.n887 Y2.n886 0.00237961
R12711 Y2.n896 Y2.n219 0.00237961
R12712 Y2.n897 Y2.n896 0.00237961
R12713 Y2.n905 Y2.n215 0.00237961
R12714 Y2.n905 Y2.n213 0.00237961
R12715 Y2.n917 Y2.n209 0.00237961
R12716 Y2.n917 Y2.n207 0.00237961
R12717 Y2.n926 Y2.n925 0.00237961
R12718 Y2.n927 Y2.n926 0.00237961
R12719 Y2.n934 Y2.n203 0.00237961
R12720 Y2.n933 Y2.n932 0.00237961
R12721 Y2.n956 Y2.n955 0.00237961
R12722 Y2.n962 Y2.n183 0.00237961
R12723 Y2.n968 Y2.n183 0.00237961
R12724 Y2.n974 Y2.n973 0.00237961
R12725 Y2.n974 Y2.n179 0.00237961
R12726 Y2.n978 Y2.n179 0.00237961
R12727 Y2.n992 Y2.n177 0.00237961
R12728 Y2.n1004 Y2.n1003 0.00237961
R12729 Y2.n1004 Y2.n167 0.00237961
R12730 Y2.n1010 Y2.n165 0.00237961
R12731 Y2.n1014 Y2.n165 0.00237961
R12732 Y2.n1014 Y2.n163 0.00237961
R12733 Y2.n1024 Y2.n1023 0.00237961
R12734 Y2.n1025 Y2.n1024 0.00237961
R12735 Y2.n1030 Y2.n159 0.00237961
R12736 Y2.n1030 Y2.n1029 0.00237961
R12737 Y2.n1059 Y2.n1058 0.00237961
R12738 Y2.n1067 Y2.n141 0.00237961
R12739 Y2.n1075 Y2.n136 0.00237961
R12740 Y2.n1080 Y2.n137 0.00237961
R12741 Y2.n1089 Y2.n132 0.00237961
R12742 Y2.n1098 Y2.n125 0.00237961
R12743 Y2.n1103 Y2.n125 0.00237961
R12744 Y2.n1108 Y2.n123 0.00237961
R12745 Y2.n1109 Y2.n1108 0.00237961
R12746 Y2.n1110 Y2.n1109 0.00237961
R12747 Y2.n1134 Y2.n121 0.00237961
R12748 Y2.n1134 Y2.n1133 0.00237961
R12749 Y2.n1128 Y2.n1127 0.00237961
R12750 Y2.n1127 Y2.n1119 0.00237961
R12751 Y2.n1151 Y2.n1150 0.00237961
R12752 Y2.n834 Y2.n248 0.00237961
R12753 Y2.n825 Y2.n264 0.00237961
R12754 Y2.n801 Y2.n298 0.00237961
R12755 Y2.n801 Y2.n800 0.00237961
R12756 Y2.n776 Y2.n775 0.00237961
R12757 Y2.n761 Y2.n760 0.00237961
R12758 Y2.n737 Y2.n398 0.00237961
R12759 Y2.n737 Y2.n736 0.00237961
R12760 Y2.n1206 Y2.n82 0.00237961
R12761 Y2.n1213 Y2.n1206 0.00237961
R12762 Y2.n1298 Y2.n1294 0.00237961
R12763 Y2.n1298 Y2.n1297 0.00237961
R12764 Y2.n953 Y2.n952 0.00235952
R12765 Y2.n965 Y2.n180 0.00235952
R12766 Y2.n253 Y2.n246 0.00235749
R12767 Y2.n854 Y2.n236 0.00235749
R12768 Y2.n866 Y2.n233 0.00235749
R12769 Y2.n874 Y2.n229 0.00235749
R12770 Y2.n882 Y2.n223 0.00235749
R12771 Y2.n909 Y2.n213 0.00235749
R12772 Y2.n934 Y2.n933 0.00235749
R12773 Y2.n955 Y2.n188 0.00235749
R12774 Y2.n962 Y2.n961 0.00235749
R12775 Y2.n992 Y2.n176 0.00235749
R12776 Y2.n1003 Y2.n169 0.00235749
R12777 Y2.n1029 Y2.n149 0.00235749
R12778 Y2.n1058 Y2.n1057 0.00235749
R12779 Y2.n1067 Y2.n143 0.00235749
R12780 Y2.n1080 Y2.n136 0.00235749
R12781 Y2.n1089 Y2.n131 0.00235749
R12782 Y2.n1098 Y2.n127 0.00235749
R12783 Y2.n1123 Y2.n1119 0.00235749
R12784 Y2.n292 Y2.n291 0.00235749
R12785 Y2.n392 Y2.n391 0.00235749
R12786 Y2.n1027 Y2.n1026 0.00233333
R12787 Y2.n909 Y2.n211 0.00231327
R12788 Y2.n1075 Y2.n139 0.00231327
R12789 Y2.n254 Y2.n251 0.00230714
R12790 Y2.n1124 Y2.n1121 0.00230714
R12791 Y2.n1120 Y2.n111 0.00230714
R12792 Y2.n927 Y2.n202 0.00229115
R12793 Y2.n1057 Y2.n147 0.00229115
R12794 Y2.n564 Y2.n533 0.00229115
R12795 Y2.n640 Y2.n639 0.00229115
R12796 Y2.n250 Y2.n237 0.00228095
R12797 Y2.n864 Y2.n230 0.00228095
R12798 Y2.n1137 Y2.n1136 0.00225476
R12799 Y2.n1053 Y2.n149 0.00224693
R12800 Y2.n820 Y2.n268 0.00222973
R12801 Y2.n756 Y2.n368 0.00222973
R12802 Y2.n100 Y2.n97 0.00222973
R12803 Y2.n1269 Y2.n1268 0.00222973
R12804 Y2.n938 Y2.n203 0.00222482
R12805 Y2.n1071 Y2.n141 0.00222482
R12806 Y2.n913 Y2.n209 0.0022027
R12807 Y2.n967 Y2.n966 0.00220238
R12808 Y2.n1011 Y2.n166 0.00220238
R12809 Y2.n983 Y2.n982 0.00217619
R12810 Y2.n990 Y2.n989 0.00217619
R12811 Y2.n877 Y2.n225 0.00215848
R12812 Y2.n1104 Y2.n123 0.00215848
R12813 Y2.n897 Y2.n217 0.00213636
R12814 Y2.n1084 Y2.n131 0.00213636
R12815 Y2.n578 Y2.n528 0.00213636
R12816 Y2.n621 Y2.n620 0.00213636
R12817 Y2.n788 Y2.n787 0.00211425
R12818 Y2.n724 Y2.n723 0.00211425
R12819 Y2.n1231 Y2.n1230 0.00211425
R12820 Y2.n1314 Y2.n48 0.00211425
R12821 Y2.n1167 Y2.n104 0.00209762
R12822 Y2.n863 Y2.n862 0.00209762
R12823 Y2.n1008 Y2.n167 0.00209214
R12824 Y2.n293 Y2.n290 0.00209214
R12825 Y2.n393 Y2.n390 0.00209214
R12826 Y2.n1189 Y2.n88 0.00209214
R12827 Y2.n1280 Y2.n1276 0.00209214
R12828 Y2.n1131 Y2.n1113 0.00207143
R12829 Y2.n951 Y2.n188 0.00207002
R12830 Y2.n973 Y2.n181 0.00207002
R12831 Y2.n1025 Y2.n158 0.00204791
R12832 Y2.n253 Y2.n252 0.0020258
R12833 Y2.n1123 Y2.n1122 0.0020258
R12834 Y2.n1150 Y2.n112 0.0020258
R12835 Y2.n958 Y2.n187 0.00201905
R12836 Y2.n808 Y2.n807 0.00201351
R12837 Y2.n744 Y2.n743 0.00201351
R12838 Y2.n1194 Y2.n87 0.00201351
R12839 Y2.n54 Y2.n14 0.00201351
R12840 Y2.n853 Y2.n238 0.00200369
R12841 Y2.n234 Y2.n231 0.00200369
R12842 Y2.n544 Y2.n537 0.00200369
R12843 Y2.n653 Y2.n509 0.00200369
R12844 Y2.n833 Y2.n260 0.00200107
R12845 Y2.n832 Y2.n831 0.00200107
R12846 Y2.n1157 Y2.n1156 0.00200107
R12847 Y2.n1022 Y2.n1021 0.00199286
R12848 Y2.n1138 Y2.n121 0.00198157
R12849 Y2.n968 Y2.n184 0.00193735
R12850 Y2.n1010 Y2.n1009 0.00193735
R12851 Y2.n981 Y2.n176 0.00191523
R12852 Y2.n988 Y2.n177 0.00191523
R12853 Y2.n834 Y2.n247 0.00191523
R12854 Y2.n830 Y2.n248 0.00191523
R12855 Y2.n1155 Y2.n107 0.00191523
R12856 Y2.n1334 Y2.n39 0.00191523
R12857 Y2.n891 Y2.n890 0.00191429
R12858 Y2.n1087 Y2.n128 0.00191429
R12859 Y2.n902 Y2.n901 0.00187101
R12860 Y2.n291 Y2.n286 0.00185493
R12861 Y2.n391 Y2.n386 0.00185493
R12862 Y2.n861 Y2.n233 0.00184889
R12863 Y2.n1083 Y2.n134 0.00184889
R12864 Y2.n597 Y2.n596 0.00184889
R12865 Y2.n605 Y2.n521 0.00184889
R12866 Y2.n827 Y2.n826 0.00184889
R12867 Y2.n356 Y2.n347 0.00184889
R12868 Y2.n762 Y2.n362 0.00184889
R12869 Y2.n459 Y2.n450 0.00184889
R12870 Y2.n1166 Y2.n1165 0.00184889
R12871 Y2.n1248 Y2.n61 0.00184889
R12872 Y2.n1263 Y2.n1259 0.00184889
R12873 Y2.n1330 Y2.n1329 0.00184889
R12874 Y2.n1062 Y2.n142 0.00183571
R12875 Y2.n1133 Y2.n1132 0.00182678
R12876 Y2.n922 Y2.n206 0.00180952
R12877 Y2.n918 Y2.n208 0.0017973
R12878 Y2.n1066 Y2.n140 0.0017973
R12879 Y2.n569 Y2.n479 0.0017973
R12880 Y2.n631 Y2.n495 0.0017973
R12881 Y2.n823 Y2.n264 0.0017897
R12882 Y2.n760 Y2.n759 0.0017897
R12883 Y2.n950 Y2.n191 0.00178256
R12884 Y2.n957 Y2.n956 0.00178256
R12885 Y2.n1035 Y2.n1034 0.00178256
R12886 Y2.n1023 Y2.n161 0.00176044
R12887 Y2.n713 Y2.n712 0.00175714
R12888 Y2.n924 Y2.n923 0.00173095
R12889 Y2.n1061 Y2.n1060 0.00173095
R12890 Y2.n870 Y2.n869 0.00171622
R12891 Y2.n775 Y2.n774 0.00171347
R12892 Y2.n892 Y2.n219 0.0016941
R12893 Y2.n132 Y2.n129 0.0016941
R12894 Y2.n1139 Y2.n120 0.0016941
R12895 Y2.n696 Y2.n695 0.0016941
R12896 Y2.n1341 Y2.n1340 0.0016941
R12897 Y2.n1095 Y2.n1094 0.00165238
R12898 Y2.n980 Y2.n979 0.00162776
R12899 Y2.n987 Y2.n986 0.00162776
R12900 Y2.n1063 Y2.n143 0.00162776
R12901 Y2.n1161 Y2.n105 0.00162776
R12902 Y2.n889 Y2.n888 0.00162619
R12903 Y2.n921 Y2.n207 0.00160565
R12904 Y2.n819 Y2.n265 0.00158354
R12905 Y2.n755 Y2.n366 0.00158354
R12906 Y2.n1172 Y2.n103 0.00158354
R12907 Y2.n1267 Y2.n1266 0.00158354
R12908 Y2.n860 Y2.n859 0.00156143
R12909 Y2.n1129 Y2.n1114 0.00156143
R12910 Y2.n588 Y2.n525 0.00156143
R12911 Y2.n612 Y2.n520 0.00156143
R12912 Y2.n777 Y2.n342 0.00156143
R12913 Y2.n711 Y2.n440 0.00156143
R12914 Y2.n1245 Y2.n1244 0.00156143
R12915 Y2.n1323 Y2.n1322 0.00156143
R12916 Y2.n959 Y2.n185 0.00154762
R12917 Y2.n1020 Y2.n162 0.00154762
R12918 Y2.n925 Y2.n205 0.00153931
R12919 Y2.n1059 Y2.n145 0.00153931
R12920 Y2.n960 Y2.n186 0.00149509
R12921 Y2.n716 Y2.n715 0.00149509
R12922 Y2.n1019 Y2.n1018 0.00147297
R12923 Y2.n1093 Y2.n127 0.00147297
R12924 Y2.n857 Y2.n235 0.00146905
R12925 Y2.n1130 Y2.n1115 0.00146905
R12926 Y2.n887 Y2.n221 0.00145086
R12927 Y2.n893 Y2.n221 0.00140663
R12928 Y2.n1093 Y2.n1092 0.00140663
R12929 Y2.n551 Y2.n534 0.00140663
R12930 Y2.n650 Y2.n649 0.00140663
R12931 Y2.n985 Y2.n984 0.00139048
R12932 Y2.n961 Y2.n960 0.00138452
R12933 Y2.n1019 Y2.n163 0.00138452
R12934 Y2.n251 Y2.n250 0.00136429
R12935 Y2.n966 Y2.n965 0.00136429
R12936 Y2.n977 Y2.n178 0.00136429
R12937 Y2.n920 Y2.n205 0.00134029
R12938 Y2.n1064 Y2.n145 0.00134029
R12939 Y2.n1007 Y2.n166 0.00133809
R12940 Y2.n1121 Y2.n1120 0.00133809
R12941 Y2.n859 Y2.n858 0.00131818
R12942 Y2.n1129 Y2.n1128 0.00131818
R12943 Y2.n777 Y2.n776 0.00131818
R12944 Y2.n1196 Y2.n86 0.00129607
R12945 Y2.n1227 Y2.n75 0.00129607
R12946 Y2.n1284 Y2.n1283 0.00129607
R12947 Y2.n1307 Y2.n49 0.00129607
R12948 Y2.n872 Y2.n871 0.00128571
R12949 Y2.n1112 Y2.n1111 0.00128571
R12950 Y2.n921 Y2.n920 0.00125184
R12951 Y2.n986 Y2.n169 0.00125184
R12952 Y2.n1064 Y2.n1063 0.00125184
R12953 Y2.n573 Y2.n572 0.00125184
R12954 Y2.n628 Y2.n627 0.00125184
R12955 Y2.n252 Y2.n238 0.00122973
R12956 Y2.n184 Y2.n181 0.00122973
R12957 Y2.n979 Y2.n978 0.00122973
R12958 Y2.n1009 Y2.n1008 0.00120762
R12959 Y2.n1122 Y2.n112 0.00120762
R12960 Y2.n931 Y2.n190 0.00120714
R12961 Y2.n1033 Y2.n1032 0.00120714
R12962 Y2.n893 Y2.n892 0.0011855
R12963 Y2.n1092 Y2.n129 0.0011855
R12964 Y2.n870 Y2.n229 0.00116339
R12965 Y2.n1110 Y2.n120 0.00116339
R12966 Y2.n816 Y2.n270 0.00114865
R12967 Y2.n752 Y2.n370 0.00114865
R12968 Y2.n1186 Y2.n91 0.00114865
R12969 Y2.n1271 Y2.n12 0.00114865
R12970 Y2.n1078 Y2.n133 0.00112857
R12971 Y2.n1018 Y2.n161 0.00111916
R12972 Y2.n900 Y2.n214 0.00110238
R12973 Y2.n932 Y2.n191 0.00109705
R12974 Y2.n957 Y2.n186 0.00109705
R12975 Y2.n1034 Y2.n159 0.00109705
R12976 Y2.n568 Y2.n567 0.00109705
R12977 Y2.n636 Y2.n632 0.00109705
R12978 Y2.n716 Y2.n439 0.00109705
R12979 Y2.n1211 Y2.n1210 0.00105283
R12980 Y2.n1303 Y2.n1302 0.00105283
R12981 Y2.n1337 Y2.n39 0.00105283
R12982 Y2.n994 Y2.n174 0.00104054
R12983 Y2.n594 Y2.n486 0.00104054
R12984 Y2.n861 Y2.n860 0.00103071
R12985 Y2.n137 Y2.n134 0.00103071
R12986 Y2.n1132 Y2.n1114 0.00103071
R12987 Y2.n258 Y2.n247 0.00103071
R12988 Y2.n826 Y2.n825 0.00103071
R12989 Y2.n762 Y2.n761 0.00103071
R12990 Y2.n1155 Y2.n109 0.00103071
R12991 Y2.n1203 Y2.n84 0.00103071
R12992 Y2.n1290 Y2.n1289 0.00103071
R12993 Y2.n901 Y2.n215 0.0010086
R12994 Y2.n981 Y2.n980 0.000964373
R12995 Y2.n988 Y2.n987 0.000964373
R12996 Y2.n830 Y2.n829 0.000964373
R12997 Y2.n461 Y2.n460 0.000964373
R12998 Y2.n1161 Y2.n1160 0.000964373
R12999 Y2.n556 Y2.n555 0.00094226
R13000 Y2.n641 Y2.n511 0.00094226
R13001 Y2.n811 Y2.n274 0.000932432
R13002 Y2.n747 Y2.n373 0.000932432
R13003 Y2.n1190 Y2.n89 0.000932432
R13004 Y2.n1277 Y2.n13 0.000932432
R13005 Y2.n834 Y2.n246 0.000898034
R13006 Y2.n1139 Y2.n1138 0.000898034
R13007 Y2.n869 Y2.n231 0.000875921
R13008 Y2.n1151 Y2.n107 0.000853808
R13009 Y2.n442 Y2.n429 0.000831695
R13010 Y2.n445 Y2.n444 0.000814286
R13011 Y2.n951 Y2.n950 0.000809582
R13012 Y2.n1035 Y2.n158 0.000809582
R13013 Y2.n581 Y2.n526 0.000787469
R13014 Y2.n617 Y2.n616 0.000787469
R13015 Y2.n293 Y2.n292 0.000787469
R13016 Y2.n393 Y2.n392 0.000787469
R13017 Y2.n443 Y2.n441 0.000765356
R13018 Y2.n99 Y2.n90 0.000765356
R13019 Y2.n1233 Y2.n1232 0.000765356
R13020 Y2.n1273 Y2.n1272 0.000765356
R13021 Y2.n1319 Y2.n1318 0.000765356
R13022 Y2.n1084 Y2.n1083 0.000743243
R13023 Y2.n902 Y2.n217 0.00072113
R13024 Y2.n868 Y2.n228 0.000716216
R13025 Y2.n1141 Y2.n1140 0.000716216
R13026 Y2.n542 Y2.n538 0.000716216
R13027 Y2.n507 Y2.n504 0.000716216
R13028 Y2.n913 Y2.n912 0.000676904
R13029 Y2.n1072 Y2.n1071 0.000654791
R13030 Y2.n540 Y2.n539 0.000654791
R13031 Y2.n505 Y2.n503 0.000654791
R13032 Y2.n1052 Y2.n147 0.000588452
R13033 Y2.n939 Y2.n202 0.000566339
R13034 Y2.n883 Y2.n882 0.000522113
R13035 Y2.n702 Y2.n458 0.000522113
R13036 nEN nEN.n1375 28.2972
R13037 nEN.n2 nEN.n1 25.6786
R13038 nEN.n1375 nEN.n2 12.7026
R13039 nEN nEN.n0 7.56318
R13040 nEN.n917 nEN.n916 2.2505
R13041 nEN.n896 nEN.n895 2.2505
R13042 nEN.n891 nEN.n337 2.2505
R13043 nEN.n889 nEN.n339 2.2505
R13044 nEN.n885 nEN.n342 2.2505
R13045 nEN.n883 nEN.n344 2.2505
R13046 nEN.n879 nEN.n347 2.2505
R13047 nEN.n877 nEN.n349 2.2505
R13048 nEN.n422 nEN.n350 2.2505
R13049 nEN.n872 nEN.n353 2.2505
R13050 nEN.n625 nEN.n355 2.2505
R13051 nEN.n866 nEN.n358 2.2505
R13052 nEN.n672 nEN.n360 2.2505
R13053 nEN.n860 nEN.n363 2.2505
R13054 nEN.n710 nEN.n365 2.2505
R13055 nEN.n1303 nEN.n1302 2.2505
R13056 nEN.n1299 nEN.n1298 2.2505
R13057 nEN.n1278 nEN.n1277 2.2505
R13058 nEN.n1275 nEN.n1274 2.2505
R13059 nEN.n1249 nEN.n1248 2.2505
R13060 nEN.n1246 nEN.n1245 2.2505
R13061 nEN.n1229 nEN.n1228 2.2505
R13062 nEN.n1227 nEN.n131 2.2505
R13063 nEN.n133 nEN.n132 2.2505
R13064 nEN.n1199 nEN.n142 2.2505
R13065 nEN.n144 nEN.n143 2.2505
R13066 nEN.n1174 nEN.n155 2.2505
R13067 nEN.n157 nEN.n156 2.2505
R13068 nEN.n1154 nEN.n167 2.2505
R13069 nEN.n169 nEN.n168 2.2505
R13070 nEN.n1304 nEN.n1303 2.2505
R13071 nEN.n1298 nEN.n1297 2.2505
R13072 nEN.n1279 nEN.n1278 2.2505
R13073 nEN.n1274 nEN.n1273 2.2505
R13074 nEN.n1250 nEN.n1249 2.2505
R13075 nEN.n1245 nEN.n1244 2.2505
R13076 nEN.n1230 nEN.n1229 2.2505
R13077 nEN.n1218 nEN.n131 2.2505
R13078 nEN.n1209 nEN.n133 2.2505
R13079 nEN.n146 nEN.n142 2.2505
R13080 nEN.n1185 nEN.n144 2.2505
R13081 nEN.n159 nEN.n155 2.2505
R13082 nEN.n1160 nEN.n157 2.2505
R13083 nEN.n177 nEN.n167 2.2505
R13084 nEN.n1141 nEN.n169 2.2505
R13085 nEN.n923 nEN.n922 2.2505
R13086 nEN.n297 nEN.n289 2.2505
R13087 nEN.n935 nEN.n285 2.2505
R13088 nEN.n944 nEN.n943 2.2505
R13089 nEN.n287 nEN.n283 2.2505
R13090 nEN.n949 nEN.n948 2.2505
R13091 nEN.n959 nEN.n271 2.2505
R13092 nEN.n968 nEN.n967 2.2505
R13093 nEN.n268 nEN.n264 2.2505
R13094 nEN.n980 nEN.n979 2.2505
R13095 nEN.n269 nEN.n257 2.2505
R13096 nEN.n975 nEN.n255 2.2505
R13097 nEN.n974 nEN.n253 2.2505
R13098 nEN.n973 nEN.n251 2.2505
R13099 nEN.n1006 nEN.n242 2.2505
R13100 nEN.n1024 nEN.n1023 2.2505
R13101 nEN.n1016 nEN.n240 2.2505
R13102 nEN.n1029 nEN.n1028 2.2505
R13103 nEN.n1032 nEN.n229 2.2505
R13104 nEN.n1048 nEN.n1047 2.2505
R13105 nEN.n231 nEN.n227 2.2505
R13106 nEN.n1053 nEN.n1052 2.2505
R13107 nEN.n1057 nEN.n216 2.2505
R13108 nEN.n1074 nEN.n1073 2.2505
R13109 nEN.n1065 nEN.n214 2.2505
R13110 nEN.n1079 nEN.n1078 2.2505
R13111 nEN.n1082 nEN.n203 2.2505
R13112 nEN.n1100 nEN.n1099 2.2505
R13113 nEN.n1092 nEN.n200 2.2505
R13114 nEN.n1106 nEN.n1105 2.2505
R13115 nEN.n201 nEN.n195 2.2505
R13116 nEN.n1120 nEN.n187 2.2505
R13117 nEN.n1134 nEN.n1133 2.2505
R13118 nEN.n185 nEN.n182 2.2505
R13119 nEN.n1136 nEN.n185 2.2505
R13120 nEN.n1135 nEN.n1134 2.2505
R13121 nEN.n187 nEN.n186 2.2505
R13122 nEN.n1103 nEN.n201 2.2505
R13123 nEN.n1105 nEN.n1104 2.2505
R13124 nEN.n1102 nEN.n200 2.2505
R13125 nEN.n1101 nEN.n1100 2.2505
R13126 nEN.n203 nEN.n202 2.2505
R13127 nEN.n1078 nEN.n1077 2.2505
R13128 nEN.n1076 nEN.n214 2.2505
R13129 nEN.n1075 nEN.n1074 2.2505
R13130 nEN.n216 nEN.n215 2.2505
R13131 nEN.n1052 nEN.n1051 2.2505
R13132 nEN.n1050 nEN.n227 2.2505
R13133 nEN.n1049 nEN.n1048 2.2505
R13134 nEN.n229 nEN.n228 2.2505
R13135 nEN.n1028 nEN.n1027 2.2505
R13136 nEN.n1026 nEN.n240 2.2505
R13137 nEN.n1025 nEN.n1024 2.2505
R13138 nEN.n242 nEN.n241 2.2505
R13139 nEN.n973 nEN.n972 2.2505
R13140 nEN.n974 nEN.n971 2.2505
R13141 nEN.n976 nEN.n975 2.2505
R13142 nEN.n977 nEN.n269 2.2505
R13143 nEN.n979 nEN.n978 2.2505
R13144 nEN.n970 nEN.n268 2.2505
R13145 nEN.n969 nEN.n968 2.2505
R13146 nEN.n271 nEN.n270 2.2505
R13147 nEN.n948 nEN.n947 2.2505
R13148 nEN.n946 nEN.n283 2.2505
R13149 nEN.n945 nEN.n944 2.2505
R13150 nEN.n285 nEN.n284 2.2505
R13151 nEN.n920 nEN.n297 2.2505
R13152 nEN.n922 nEN.n921 2.2505
R13153 nEN.n918 nEN.n917 2.2505
R13154 nEN.n895 nEN.n894 2.2505
R13155 nEN.n892 nEN.n891 2.2505
R13156 nEN.n889 nEN.n888 2.2505
R13157 nEN.n886 nEN.n885 2.2505
R13158 nEN.n883 nEN.n882 2.2505
R13159 nEN.n880 nEN.n879 2.2505
R13160 nEN.n877 nEN.n876 2.2505
R13161 nEN.n875 nEN.n350 2.2505
R13162 nEN.n872 nEN.n351 2.2505
R13163 nEN.n869 nEN.n355 2.2505
R13164 nEN.n866 nEN.n356 2.2505
R13165 nEN.n863 nEN.n360 2.2505
R13166 nEN.n860 nEN.n361 2.2505
R13167 nEN.n857 nEN.n365 2.2505
R13168 nEN.n1316 nEN.n86 2.2505
R13169 nEN.n1317 nEN.n85 2.2505
R13170 nEN.n84 nEN.n82 2.2505
R13171 nEN.n83 nEN.n67 2.2505
R13172 nEN.n1329 nEN.n66 2.2505
R13173 nEN.n1330 nEN.n65 2.2505
R13174 nEN.n64 nEN.n62 2.2505
R13175 nEN.n63 nEN.n40 2.2505
R13176 nEN.n1342 nEN.n39 2.2505
R13177 nEN.n1343 nEN.n38 2.2505
R13178 nEN.n37 nEN.n33 2.2505
R13179 nEN.n36 nEN.n35 2.2505
R13180 nEN.n34 nEN.n22 2.2505
R13181 nEN.n1359 nEN.n21 2.2505
R13182 nEN.n1360 nEN.n20 2.2505
R13183 nEN.n19 nEN.n7 2.2505
R13184 nEN.n1371 nEN.n3 2.2505
R13185 nEN.n791 nEN.n4 2.2505
R13186 nEN.n778 nEN.n777 2.2505
R13187 nEN.n811 nEN.n776 2.2505
R13188 nEN.n812 nEN.n775 2.2505
R13189 nEN.n774 nEN.n772 2.2505
R13190 nEN.n773 nEN.n750 2.2505
R13191 nEN.n824 nEN.n749 2.2505
R13192 nEN.n825 nEN.n748 2.2505
R13193 nEN.n747 nEN.n743 2.2505
R13194 nEN.n746 nEN.n745 2.2505
R13195 nEN.n744 nEN.n732 2.2505
R13196 nEN.n841 nEN.n731 2.2505
R13197 nEN.n842 nEN.n730 2.2505
R13198 nEN.n729 nEN.n368 2.2505
R13199 nEN.n854 nEN.n366 2.2505
R13200 nEN.n854 nEN.n853 2.2505
R13201 nEN.n726 nEN.n368 2.2505
R13202 nEN.n843 nEN.n842 2.2505
R13203 nEN.n841 nEN.n840 2.2505
R13204 nEN.n734 nEN.n732 2.2505
R13205 nEN.n745 nEN.n738 2.2505
R13206 nEN.n743 nEN.n740 2.2505
R13207 nEN.n826 nEN.n825 2.2505
R13208 nEN.n824 nEN.n823 2.2505
R13209 nEN.n767 nEN.n750 2.2505
R13210 nEN.n772 nEN.n771 2.2505
R13211 nEN.n813 nEN.n812 2.2505
R13212 nEN.n811 nEN.n810 2.2505
R13213 nEN.n787 nEN.n778 2.2505
R13214 nEN.n792 nEN.n791 2.2505
R13215 nEN.n800 nEN.n5 2.2505
R13216 nEN.n1372 nEN.n6 2.2505
R13217 nEN.n1371 nEN.n1370 2.2505
R13218 nEN.n16 nEN.n7 2.2505
R13219 nEN.n1361 nEN.n1360 2.2505
R13220 nEN.n1359 nEN.n1358 2.2505
R13221 nEN.n24 nEN.n22 2.2505
R13222 nEN.n35 nEN.n28 2.2505
R13223 nEN.n33 nEN.n30 2.2505
R13224 nEN.n1344 nEN.n1343 2.2505
R13225 nEN.n1342 nEN.n1341 2.2505
R13226 nEN.n57 nEN.n40 2.2505
R13227 nEN.n62 nEN.n61 2.2505
R13228 nEN.n1331 nEN.n1330 2.2505
R13229 nEN.n1329 nEN.n1328 2.2505
R13230 nEN.n76 nEN.n67 2.2505
R13231 nEN.n82 nEN.n80 2.2505
R13232 nEN.n1318 nEN.n1317 2.2505
R13233 nEN.n1316 nEN.n1315 2.2505
R13234 nEN.n712 nEN.n711 2.2005
R13235 nEN.n709 nEN.n708 2.2005
R13236 nEN.n703 nEN.n382 2.2005
R13237 nEN.n389 nEN.n386 2.2005
R13238 nEN.n696 nEN.n390 2.2005
R13239 nEN.n691 nEN.n690 2.2005
R13240 nEN.n681 nEN.n392 2.2005
R13241 nEN.n683 nEN.n682 2.2005
R13242 nEN.n673 nEN.n394 2.2005
R13243 nEN.n675 nEN.n674 2.2005
R13244 nEN.n671 nEN.n670 2.2005
R13245 nEN.n663 nEN.n397 2.2005
R13246 nEN.n657 nEN.n656 2.2005
R13247 nEN.n655 nEN.n654 2.2005
R13248 nEN.n650 nEN.n649 2.2005
R13249 nEN.n648 nEN.n647 2.2005
R13250 nEN.n642 nEN.n641 2.2005
R13251 nEN.n640 nEN.n639 2.2005
R13252 nEN.n633 nEN.n409 2.2005
R13253 nEN.n627 nEN.n626 2.2005
R13254 nEN.n624 nEN.n623 2.2005
R13255 nEN.n614 nEN.n414 2.2005
R13256 nEN.n616 nEN.n615 2.2005
R13257 nEN.n609 nEN.n608 2.2005
R13258 nEN.n607 nEN.n606 2.2005
R13259 nEN.n600 nEN.n599 2.2005
R13260 nEN.n598 nEN.n597 2.2005
R13261 nEN.n591 nEN.n590 2.2005
R13262 nEN.n589 nEN.n588 2.2005
R13263 nEN.n582 nEN.n581 2.2005
R13264 nEN.n580 nEN.n579 2.2005
R13265 nEN.n573 nEN.n572 2.2005
R13266 nEN.n571 nEN.n570 2.2005
R13267 nEN.n565 nEN.n433 2.2005
R13268 nEN.n556 nEN.n437 2.2005
R13269 nEN.n558 nEN.n557 2.2005
R13270 nEN.n554 nEN.n553 2.2005
R13271 nEN.n546 nEN.n440 2.2005
R13272 nEN.n540 nEN.n539 2.2005
R13273 nEN.n538 nEN.n537 2.2005
R13274 nEN.n533 nEN.n532 2.2005
R13275 nEN.n531 nEN.n530 2.2005
R13276 nEN.n525 nEN.n524 2.2005
R13277 nEN.n523 nEN.n522 2.2005
R13278 nEN.n516 nEN.n452 2.2005
R13279 nEN.n510 nEN.n509 2.2005
R13280 nEN.n507 nEN.n506 2.2005
R13281 nEN.n497 nEN.n457 2.2005
R13282 nEN.n499 nEN.n498 2.2005
R13283 nEN.n492 nEN.n491 2.2005
R13284 nEN.n490 nEN.n489 2.2005
R13285 nEN.n483 nEN.n482 2.2005
R13286 nEN.n481 nEN.n480 2.2005
R13287 nEN.n474 nEN.n473 2.2005
R13288 nEN.n471 nEN.n334 2.2005
R13289 nEN.n898 nEN.n897 2.2005
R13290 nEN.n903 nEN.n330 2.2005
R13291 nEN.n329 nEN.n326 2.2005
R13292 nEN.n910 nEN.n301 2.2005
R13293 nEN.n915 nEN.n914 2.2005
R13294 nEN.n321 nEN.n300 2.2005
R13295 nEN.n90 nEN.n89 2.2005
R13296 nEN.n1140 nEN.n181 2.2005
R13297 nEN.n1143 nEN.n1142 2.2005
R13298 nEN.n172 nEN.n170 2.2005
R13299 nEN.n1150 nEN.n1149 2.2005
R13300 nEN.n1148 nEN.n171 2.2005
R13301 nEN.n179 nEN.n178 2.2005
R13302 nEN.n176 nEN.n175 2.2005
R13303 nEN.n173 nEN.n166 2.2005
R13304 nEN.n1158 nEN.n163 2.2005
R13305 nEN.n1162 nEN.n1161 2.2005
R13306 nEN.n1159 nEN.n165 2.2005
R13307 nEN.n164 nEN.n158 2.2005
R13308 nEN.n1170 nEN.n1169 2.2005
R13309 nEN.n1168 nEN.n160 2.2005
R13310 nEN.n154 nEN.n153 2.2005
R13311 nEN.n1179 nEN.n1178 2.2005
R13312 nEN.n1181 nEN.n152 2.2005
R13313 nEN.n1183 nEN.n1182 2.2005
R13314 nEN.n1184 nEN.n150 2.2005
R13315 nEN.n1187 nEN.n1186 2.2005
R13316 nEN.n151 nEN.n145 2.2005
R13317 nEN.n1195 nEN.n1194 2.2005
R13318 nEN.n1193 nEN.n147 2.2005
R13319 nEN.n141 nEN.n140 2.2005
R13320 nEN.n1204 nEN.n1203 2.2005
R13321 nEN.n1205 nEN.n139 2.2005
R13322 nEN.n1208 nEN.n1207 2.2005
R13323 nEN.n1210 nEN.n138 2.2005
R13324 nEN.n1212 nEN.n1211 2.2005
R13325 nEN.n136 nEN.n134 2.2005
R13326 nEN.n1223 nEN.n1222 2.2005
R13327 nEN.n1221 nEN.n135 2.2005
R13328 nEN.n1220 nEN.n1219 2.2005
R13329 nEN.n1216 nEN.n130 2.2005
R13330 nEN.n1231 nEN.n127 2.2005
R13331 nEN.n1235 nEN.n1234 2.2005
R13332 nEN.n1232 nEN.n129 2.2005
R13333 nEN.n128 nEN.n122 2.2005
R13334 nEN.n1243 nEN.n1242 2.2005
R13335 nEN.n1241 nEN.n124 2.2005
R13336 nEN.n118 nEN.n117 2.2005
R13337 nEN.n1252 nEN.n1251 2.2005
R13338 nEN.n1254 nEN.n116 2.2005
R13339 nEN.n1256 nEN.n1255 2.2005
R13340 nEN.n1257 nEN.n115 2.2005
R13341 nEN.n1260 nEN.n1259 2.2005
R13342 nEN.n113 nEN.n111 2.2005
R13343 nEN.n1272 nEN.n1271 2.2005
R13344 nEN.n1270 nEN.n112 2.2005
R13345 nEN.n1268 nEN.n1267 2.2005
R13346 nEN.n1265 nEN.n107 2.2005
R13347 nEN.n1280 nEN.n106 2.2005
R13348 nEN.n1284 nEN.n1283 2.2005
R13349 nEN.n1281 nEN.n104 2.2005
R13350 nEN.n1289 nEN.n102 2.2005
R13351 nEN.n1296 nEN.n1295 2.2005
R13352 nEN.n1293 nEN.n103 2.2005
R13353 nEN.n1292 nEN.n1291 2.2005
R13354 nEN.n98 nEN.n97 2.2005
R13355 nEN.n1306 nEN.n1305 2.2005
R13356 nEN.n373 nEN.n369 2.2005
R13357 nEN.n852 nEN.n851 2.2005
R13358 nEN.n722 nEN.n370 2.2005
R13359 nEN.n727 nEN.n724 2.2005
R13360 nEN.n845 nEN.n844 2.2005
R13361 nEN.n728 nEN.n725 2.2005
R13362 nEN.n735 nEN.n733 2.2005
R13363 nEN.n839 nEN.n838 2.2005
R13364 nEN.n837 nEN.n836 2.2005
R13365 nEN.n835 nEN.n834 2.2005
R13366 nEN.n833 nEN.n832 2.2005
R13367 nEN.n831 nEN.n830 2.2005
R13368 nEN.n829 nEN.n828 2.2005
R13369 nEN.n827 nEN.n741 2.2005
R13370 nEN.n758 nEN.n742 2.2005
R13371 nEN.n757 nEN.n751 2.2005
R13372 nEN.n822 nEN.n821 2.2005
R13373 nEN.n820 nEN.n752 2.2005
R13374 nEN.n768 nEN.n754 2.2005
R13375 nEN.n770 nEN.n769 2.2005
R13376 nEN.n765 nEN.n763 2.2005
R13377 nEN.n815 nEN.n814 2.2005
R13378 nEN.n766 nEN.n764 2.2005
R13379 nEN.n782 nEN.n779 2.2005
R13380 nEN.n809 nEN.n808 2.2005
R13381 nEN.n783 nEN.n780 2.2005
R13382 nEN.n789 nEN.n788 2.2005
R13383 nEN.n790 nEN.n785 2.2005
R13384 nEN.n803 nEN.n802 2.2005
R13385 nEN.n801 nEN.n786 2.2005
R13386 nEN.n799 nEN.n798 2.2005
R13387 nEN.n797 nEN.n793 2.2005
R13388 nEN.n796 nEN.n795 2.2005
R13389 nEN.n10 nEN.n8 2.2005
R13390 nEN.n1369 nEN.n1368 2.2005
R13391 nEN.n11 nEN.n9 2.2005
R13392 nEN.n17 nEN.n14 2.2005
R13393 nEN.n1363 nEN.n1362 2.2005
R13394 nEN.n18 nEN.n15 2.2005
R13395 nEN.n25 nEN.n23 2.2005
R13396 nEN.n1357 nEN.n1356 2.2005
R13397 nEN.n1355 nEN.n1354 2.2005
R13398 nEN.n1353 nEN.n1352 2.2005
R13399 nEN.n1351 nEN.n1350 2.2005
R13400 nEN.n1349 nEN.n1348 2.2005
R13401 nEN.n1347 nEN.n1346 2.2005
R13402 nEN.n1345 nEN.n31 2.2005
R13403 nEN.n48 nEN.n32 2.2005
R13404 nEN.n47 nEN.n41 2.2005
R13405 nEN.n1340 nEN.n1339 2.2005
R13406 nEN.n1338 nEN.n42 2.2005
R13407 nEN.n58 nEN.n44 2.2005
R13408 nEN.n60 nEN.n59 2.2005
R13409 nEN.n55 nEN.n53 2.2005
R13410 nEN.n1333 nEN.n1332 2.2005
R13411 nEN.n56 nEN.n54 2.2005
R13412 nEN.n71 nEN.n68 2.2005
R13413 nEN.n1327 nEN.n1326 2.2005
R13414 nEN.n72 nEN.n69 2.2005
R13415 nEN.n78 nEN.n77 2.2005
R13416 nEN.n79 nEN.n74 2.2005
R13417 nEN.n1321 nEN.n1320 2.2005
R13418 nEN.n1319 nEN.n75 2.2005
R13419 nEN.n92 nEN.n81 2.2005
R13420 nEN.n93 nEN.n88 2.2005
R13421 nEN.n309 nEN.n295 2.2005
R13422 nEN.n924 nEN.n294 2.2005
R13423 nEN.n926 nEN.n925 2.2005
R13424 nEN.n933 nEN.n932 2.2005
R13425 nEN.n934 nEN.n288 2.2005
R13426 nEN.n937 nEN.n936 2.2005
R13427 nEN.n939 nEN.n286 2.2005
R13428 nEN.n942 nEN.n941 2.2005
R13429 nEN.n282 nEN.n280 2.2005
R13430 nEN.n951 nEN.n950 2.2005
R13431 nEN.n276 nEN.n275 2.2005
R13432 nEN.n958 nEN.n957 2.2005
R13433 nEN.n961 nEN.n960 2.2005
R13434 nEN.n963 nEN.n272 2.2005
R13435 nEN.n966 nEN.n965 2.2005
R13436 nEN.n273 nEN.n262 2.2005
R13437 nEN.n983 nEN.n982 2.2005
R13438 nEN.n981 nEN.n263 2.2005
R13439 nEN.n267 nEN.n266 2.2005
R13440 nEN.n265 nEN.n258 2.2005
R13441 nEN.n991 nEN.n990 2.2005
R13442 nEN.n993 nEN.n992 2.2005
R13443 nEN.n995 nEN.n994 2.2005
R13444 nEN.n997 nEN.n996 2.2005
R13445 nEN.n999 nEN.n998 2.2005
R13446 nEN.n1001 nEN.n1000 2.2005
R13447 nEN.n1004 nEN.n1003 2.2005
R13448 nEN.n1005 nEN.n249 2.2005
R13449 nEN.n1008 nEN.n1007 2.2005
R13450 nEN.n245 nEN.n243 2.2005
R13451 nEN.n1022 nEN.n1021 2.2005
R13452 nEN.n1020 nEN.n244 2.2005
R13453 nEN.n1018 nEN.n1017 2.2005
R13454 nEN.n1014 nEN.n239 2.2005
R13455 nEN.n1030 nEN.n237 2.2005
R13456 nEN.n1034 nEN.n1033 2.2005
R13457 nEN.n1031 nEN.n233 2.2005
R13458 nEN.n1040 nEN.n230 2.2005
R13459 nEN.n1046 nEN.n1045 2.2005
R13460 nEN.n1043 nEN.n232 2.2005
R13461 nEN.n1041 nEN.n226 2.2005
R13462 nEN.n1054 nEN.n224 2.2005
R13463 nEN.n1059 nEN.n1058 2.2005
R13464 nEN.n1056 nEN.n1055 2.2005
R13465 nEN.n219 nEN.n217 2.2005
R13466 nEN.n1072 nEN.n1071 2.2005
R13467 nEN.n1069 nEN.n218 2.2005
R13468 nEN.n1067 nEN.n1066 2.2005
R13469 nEN.n213 nEN.n211 2.2005
R13470 nEN.n1085 nEN.n1084 2.2005
R13471 nEN.n1083 nEN.n212 2.2005
R13472 nEN.n1081 nEN.n1080 2.2005
R13473 nEN.n208 nEN.n204 2.2005
R13474 nEN.n1098 nEN.n1097 2.2005
R13475 nEN.n1095 nEN.n205 2.2005
R13476 nEN.n1094 nEN.n1093 2.2005
R13477 nEN.n199 nEN.n198 2.2005
R13478 nEN.n1109 nEN.n1108 2.2005
R13479 nEN.n1107 nEN.n196 2.2005
R13480 nEN.n1118 nEN.n1117 2.2005
R13481 nEN.n1122 nEN.n1121 2.2005
R13482 nEN.n1119 nEN.n192 2.2005
R13483 nEN.n191 nEN.n188 2.2005
R13484 nEN.n1132 nEN.n1131 2.2005
R13485 nEN.n1130 nEN.n189 2.2005
R13486 nEN.n328 nEN.n299 1.8005
R13487 nEN.n465 nEN.n335 1.8005
R13488 nEN.n890 nEN.n338 1.8005
R13489 nEN.n508 nEN.n340 1.8005
R13490 nEN.n884 nEN.n343 1.8005
R13491 nEN.n555 nEN.n345 1.8005
R13492 nEN.n878 nEN.n348 1.8005
R13493 nEN.n873 nEN.n352 1.8005
R13494 nEN.n871 nEN.n354 1.8005
R13495 nEN.n867 nEN.n357 1.8005
R13496 nEN.n865 nEN.n359 1.8005
R13497 nEN.n861 nEN.n362 1.8005
R13498 nEN.n859 nEN.n364 1.8005
R13499 nEN.n1300 nEN.n99 1.8005
R13500 nEN.n101 nEN.n100 1.8005
R13501 nEN.n1276 nEN.n108 1.8005
R13502 nEN.n110 nEN.n109 1.8005
R13503 nEN.n1247 nEN.n119 1.8005
R13504 nEN.n121 nEN.n120 1.8005
R13505 nEN.n1226 nEN.n1225 1.8005
R13506 nEN.n1201 nEN.n1200 1.8005
R13507 nEN.n1198 nEN.n1197 1.8005
R13508 nEN.n1176 nEN.n1175 1.8005
R13509 nEN.n1173 nEN.n1172 1.8005
R13510 nEN.n1156 nEN.n1155 1.8005
R13511 nEN.n1153 nEN.n1152 1.8005
R13512 nEN.n1290 nEN.n99 1.8005
R13513 nEN.n1282 nEN.n101 1.8005
R13514 nEN.n1266 nEN.n108 1.8005
R13515 nEN.n1258 nEN.n110 1.8005
R13516 nEN.n123 nEN.n119 1.8005
R13517 nEN.n1233 nEN.n121 1.8005
R13518 nEN.n1225 nEN.n1224 1.8005
R13519 nEN.n1202 nEN.n1201 1.8005
R13520 nEN.n1197 nEN.n1196 1.8005
R13521 nEN.n1177 nEN.n1176 1.8005
R13522 nEN.n1172 nEN.n1171 1.8005
R13523 nEN.n1157 nEN.n1156 1.8005
R13524 nEN.n1152 nEN.n1151 1.8005
R13525 nEN.n1139 nEN.n1138 1.8005
R13526 nEN.n1138 nEN.n1137 1.8005
R13527 nEN.n299 nEN.n298 1.8005
R13528 nEN.n893 nEN.n335 1.8005
R13529 nEN.n890 nEN.n336 1.8005
R13530 nEN.n887 nEN.n340 1.8005
R13531 nEN.n884 nEN.n341 1.8005
R13532 nEN.n881 nEN.n345 1.8005
R13533 nEN.n878 nEN.n346 1.8005
R13534 nEN.n874 nEN.n873 1.8005
R13535 nEN.n871 nEN.n870 1.8005
R13536 nEN.n868 nEN.n867 1.8005
R13537 nEN.n865 nEN.n864 1.8005
R13538 nEN.n862 nEN.n861 1.8005
R13539 nEN.n859 nEN.n858 1.8005
R13540 nEN.n1301 nEN.n87 1.8005
R13541 nEN.n1314 nEN.n87 1.8005
R13542 nEN.n305 nEN.n296 1.5005
R13543 nEN.n919 nEN.n296 1.5005
R13544 nEN.n856 nEN.n855 1.5005
R13545 nEN.n855 nEN.n367 1.5005
R13546 nEN.n1374 nEN.n1373 1.11718
R13547 nEN.n721 nEN.n371 1.1125
R13548 nEN.n1114 nEN.n194 1.10836
R13549 nEN.n1116 nEN.n1115 1.10443
R13550 nEN.n1129 nEN.n1128 1.10381
R13551 nEN.n720 nEN.n374 1.10372
R13552 nEN.n1110 nEN.n197 1.10339
R13553 nEN.n1125 nEN.n192 1.10272
R13554 nEN.n1122 nEN.n193 1.10272
R13555 nEN.n1113 nEN.n196 1.10272
R13556 nEN.n851 nEN.n850 1.10263
R13557 nEN.n848 nEN.n722 1.10263
R13558 nEN.n1308 nEN.n1307 1.1005
R13559 nEN.n1145 nEN.n1144 1.1005
R13560 nEN.n1147 nEN.n1146 1.1005
R13561 nEN.n174 nEN.n162 1.1005
R13562 nEN.n1164 nEN.n1163 1.1005
R13563 nEN.n1165 nEN.n161 1.1005
R13564 nEN.n1167 nEN.n1166 1.1005
R13565 nEN.n1180 nEN.n149 1.1005
R13566 nEN.n1189 nEN.n1188 1.1005
R13567 nEN.n1190 nEN.n148 1.1005
R13568 nEN.n1192 nEN.n1191 1.1005
R13569 nEN.n1206 nEN.n137 1.1005
R13570 nEN.n1214 nEN.n1213 1.1005
R13571 nEN.n1222 nEN.n1215 1.1005
R13572 nEN.n1217 nEN.n126 1.1005
R13573 nEN.n1237 nEN.n1236 1.1005
R13574 nEN.n1238 nEN.n125 1.1005
R13575 nEN.n1240 nEN.n1239 1.1005
R13576 nEN.n1253 nEN.n114 1.1005
R13577 nEN.n1262 nEN.n1261 1.1005
R13578 nEN.n1264 nEN.n1263 1.1005
R13579 nEN.n1269 nEN.n105 1.1005
R13580 nEN.n1286 nEN.n1285 1.1005
R13581 nEN.n1288 nEN.n1287 1.1005
R13582 nEN.n1294 nEN.n96 1.1005
R13583 nEN.n183 nEN.n180 1.1005
R13584 nEN.n95 nEN.n94 1.1005
R13585 nEN.n1311 nEN.n1310 1.1005
R13586 nEN.n1310 nEN.n1309 1.1005
R13587 nEN.n1313 nEN.n1312 1.1005
R13588 nEN.n91 nEN.n73 1.1005
R13589 nEN.n1323 nEN.n1322 1.1005
R13590 nEN.n1325 nEN.n1324 1.1005
R13591 nEN.n70 nEN.n52 1.1005
R13592 nEN.n1335 nEN.n1334 1.1005
R13593 nEN.n1337 nEN.n1336 1.1005
R13594 nEN.n51 nEN.n43 1.1005
R13595 nEN.n50 nEN.n49 1.1005
R13596 nEN.n46 nEN.n29 1.1005
R13597 nEN.n45 nEN.n27 1.1005
R13598 nEN.n26 nEN.n13 1.1005
R13599 nEN.n1365 nEN.n1364 1.1005
R13600 nEN.n1367 nEN.n1366 1.1005
R13601 nEN.n796 nEN.n12 1.1005
R13602 nEN.n794 nEN.n784 1.1005
R13603 nEN.n805 nEN.n804 1.1005
R13604 nEN.n807 nEN.n806 1.1005
R13605 nEN.n781 nEN.n762 1.1005
R13606 nEN.n817 nEN.n816 1.1005
R13607 nEN.n819 nEN.n818 1.1005
R13608 nEN.n761 nEN.n753 1.1005
R13609 nEN.n760 nEN.n759 1.1005
R13610 nEN.n756 nEN.n739 1.1005
R13611 nEN.n755 nEN.n737 1.1005
R13612 nEN.n736 nEN.n723 1.1005
R13613 nEN.n847 nEN.n846 1.1005
R13614 nEN.n849 nEN.n372 1.1005
R13615 nEN.n717 nEN.n375 1.1005
R13616 nEN.n719 nEN.n718 1.1005
R13617 nEN.n378 nEN.n377 1.1005
R13618 nEN.n717 nEN.n716 1.1005
R13619 nEN.n713 nEN.n712 1.1005
R13620 nEN.n706 nEN.n384 1.1005
R13621 nEN.n708 nEN.n707 1.1005
R13622 nEN.n704 nEN.n703 1.1005
R13623 nEN.n701 nEN.n700 1.1005
R13624 nEN.n697 nEN.n387 1.1005
R13625 nEN.n696 nEN.n695 1.1005
R13626 nEN.n694 nEN.n388 1.1005
R13627 nEN.n688 nEN.n687 1.1005
R13628 nEN.n677 nEN.n676 1.1005
R13629 nEN.n675 nEN.n395 1.1005
R13630 nEN.n667 nEN.n396 1.1005
R13631 nEN.n665 nEN.n664 1.1005
R13632 nEN.n663 nEN.n399 1.1005
R13633 nEN.n662 nEN.n661 1.1005
R13634 nEN.n402 nEN.n401 1.1005
R13635 nEN.n644 nEN.n406 1.1005
R13636 nEN.n643 nEN.n642 1.1005
R13637 nEN.n408 nEN.n407 1.1005
R13638 nEN.n635 nEN.n634 1.1005
R13639 nEN.n633 nEN.n411 1.1005
R13640 nEN.n632 nEN.n631 1.1005
R13641 nEN.n629 nEN.n628 1.1005
R13642 nEN.n623 nEN.n413 1.1005
R13643 nEN.n620 nEN.n414 1.1005
R13644 nEN.n617 nEN.n415 1.1005
R13645 nEN.n611 nEN.n416 1.1005
R13646 nEN.n610 nEN.n609 1.1005
R13647 nEN.n418 nEN.n417 1.1005
R13648 nEN.n602 nEN.n601 1.1005
R13649 nEN.n593 nEN.n592 1.1005
R13650 nEN.n591 nEN.n424 1.1005
R13651 nEN.n588 nEN.n587 1.1005
R13652 nEN.n584 nEN.n583 1.1005
R13653 nEN.n577 nEN.n430 1.1005
R13654 nEN.n579 nEN.n578 1.1005
R13655 nEN.n576 nEN.n429 1.1005
R13656 nEN.n568 nEN.n435 1.1005
R13657 nEN.n563 nEN.n562 1.1005
R13658 nEN.n561 nEN.n437 1.1005
R13659 nEN.n558 nEN.n438 1.1005
R13660 nEN.n552 nEN.n551 1.1005
R13661 nEN.n548 nEN.n547 1.1005
R13662 nEN.n546 nEN.n442 1.1005
R13663 nEN.n545 nEN.n544 1.1005
R13664 nEN.n445 nEN.n444 1.1005
R13665 nEN.n527 nEN.n449 1.1005
R13666 nEN.n526 nEN.n525 1.1005
R13667 nEN.n451 nEN.n450 1.1005
R13668 nEN.n518 nEN.n517 1.1005
R13669 nEN.n516 nEN.n454 1.1005
R13670 nEN.n515 nEN.n514 1.1005
R13671 nEN.n512 nEN.n511 1.1005
R13672 nEN.n506 nEN.n456 1.1005
R13673 nEN.n503 nEN.n457 1.1005
R13674 nEN.n500 nEN.n458 1.1005
R13675 nEN.n494 nEN.n459 1.1005
R13676 nEN.n493 nEN.n492 1.1005
R13677 nEN.n461 nEN.n460 1.1005
R13678 nEN.n485 nEN.n484 1.1005
R13679 nEN.n483 nEN.n463 1.1005
R13680 nEN.n477 nEN.n464 1.1005
R13681 nEN.n476 nEN.n466 1.1005
R13682 nEN.n475 nEN.n474 1.1005
R13683 nEN.n471 nEN.n470 1.1005
R13684 nEN.n333 nEN.n332 1.1005
R13685 nEN.n901 nEN.n331 1.1005
R13686 nEN.n903 nEN.n902 1.1005
R13687 nEN.n904 nEN.n327 1.1005
R13688 nEN.n909 nEN.n325 1.1005
R13689 nEN.n323 nEN.n322 1.1005
R13690 nEN.n321 nEN.n304 1.1005
R13691 nEN.n320 nEN.n319 1.1005
R13692 nEN.n911 nEN.n910 1.1005
R13693 nEN.n912 nEN.n303 1.1005
R13694 nEN.n914 nEN.n913 1.1005
R13695 nEN.n324 nEN.n302 1.1005
R13696 nEN.n908 nEN.n907 1.1005
R13697 nEN.n906 nEN.n905 1.1005
R13698 nEN.n900 nEN.n899 1.1005
R13699 nEN.n469 nEN.n468 1.1005
R13700 nEN.n472 nEN.n467 1.1005
R13701 nEN.n479 nEN.n478 1.1005
R13702 nEN.n486 nEN.n462 1.1005
R13703 nEN.n488 nEN.n487 1.1005
R13704 nEN.n496 nEN.n495 1.1005
R13705 nEN.n502 nEN.n501 1.1005
R13706 nEN.n505 nEN.n504 1.1005
R13707 nEN.n513 nEN.n455 1.1005
R13708 nEN.n519 nEN.n453 1.1005
R13709 nEN.n521 nEN.n520 1.1005
R13710 nEN.n529 nEN.n528 1.1005
R13711 nEN.n537 nEN.n536 1.1005
R13712 nEN.n535 nEN.n446 1.1005
R13713 nEN.n534 nEN.n533 1.1005
R13714 nEN.n448 nEN.n447 1.1005
R13715 nEN.n542 nEN.n541 1.1005
R13716 nEN.n543 nEN.n443 1.1005
R13717 nEN.n549 nEN.n441 1.1005
R13718 nEN.n550 nEN.n439 1.1005
R13719 nEN.n560 nEN.n559 1.1005
R13720 nEN.n570 nEN.n569 1.1005
R13721 nEN.n567 nEN.n434 1.1005
R13722 nEN.n566 nEN.n565 1.1005
R13723 nEN.n564 nEN.n436 1.1005
R13724 nEN.n432 nEN.n431 1.1005
R13725 nEN.n575 nEN.n574 1.1005
R13726 nEN.n428 nEN.n427 1.1005
R13727 nEN.n585 nEN.n426 1.1005
R13728 nEN.n586 nEN.n425 1.1005
R13729 nEN.n600 nEN.n420 1.1005
R13730 nEN.n595 nEN.n421 1.1005
R13731 nEN.n597 nEN.n596 1.1005
R13732 nEN.n594 nEN.n423 1.1005
R13733 nEN.n603 nEN.n419 1.1005
R13734 nEN.n605 nEN.n604 1.1005
R13735 nEN.n613 nEN.n612 1.1005
R13736 nEN.n619 nEN.n618 1.1005
R13737 nEN.n622 nEN.n621 1.1005
R13738 nEN.n630 nEN.n412 1.1005
R13739 nEN.n636 nEN.n410 1.1005
R13740 nEN.n638 nEN.n637 1.1005
R13741 nEN.n646 nEN.n645 1.1005
R13742 nEN.n654 nEN.n653 1.1005
R13743 nEN.n652 nEN.n403 1.1005
R13744 nEN.n651 nEN.n650 1.1005
R13745 nEN.n405 nEN.n404 1.1005
R13746 nEN.n659 nEN.n658 1.1005
R13747 nEN.n660 nEN.n400 1.1005
R13748 nEN.n666 nEN.n398 1.1005
R13749 nEN.n669 nEN.n668 1.1005
R13750 nEN.n678 nEN.n394 1.1005
R13751 nEN.n686 nEN.n392 1.1005
R13752 nEN.n685 nEN.n684 1.1005
R13753 nEN.n683 nEN.n393 1.1005
R13754 nEN.n680 nEN.n679 1.1005
R13755 nEN.n689 nEN.n391 1.1005
R13756 nEN.n693 nEN.n692 1.1005
R13757 nEN.n699 nEN.n698 1.1005
R13758 nEN.n702 nEN.n385 1.1005
R13759 nEN.n705 nEN.n383 1.1005
R13760 nEN.n715 nEN.n377 1.1005
R13761 nEN.n381 nEN.n380 1.1005
R13762 nEN.n714 nEN.n376 1.1005
R13763 nEN.n312 nEN.n311 1.1005
R13764 nEN.n927 nEN.n292 1.1005
R13765 nEN.n952 nEN.n278 1.1005
R13766 nEN.n1009 nEN.n247 1.1005
R13767 nEN.n1035 nEN.n235 1.1005
R13768 nEN.n1060 nEN.n222 1.1005
R13769 nEN.n308 nEN.n307 1.1005
R13770 nEN.n317 nEN.n314 1.1005
R13771 nEN.n310 nEN.n293 1.1005
R13772 nEN.n1126 nEN.n190 1.1005
R13773 nEN.n1124 nEN.n1123 1.1005
R13774 nEN.n1112 nEN.n1111 1.1005
R13775 nEN.n1091 nEN.n1090 1.1005
R13776 nEN.n1087 nEN.n1086 1.1005
R13777 nEN.n1062 nEN.n1061 1.1005
R13778 nEN.n1039 nEN.n1038 1.1005
R13779 nEN.n1037 nEN.n1036 1.1005
R13780 nEN.n1013 nEN.n1012 1.1005
R13781 nEN.n1011 nEN.n1010 1.1005
R13782 nEN.n987 nEN.n254 1.1005
R13783 nEN.n985 nEN.n984 1.1005
R13784 nEN.n954 nEN.n953 1.1005
R13785 nEN.n931 nEN.n930 1.1005
R13786 nEN.n929 nEN.n928 1.1005
R13787 nEN.n313 nEN.n306 1.1005
R13788 nEN.n315 nEN.n308 1.1005
R13789 nEN.n318 nEN.n317 1.1005
R13790 nEN.n1314 nEN.n1313 0.733833
R13791 nEN.n718 nEN.n367 0.733833
R13792 nEN.n306 nEN.n305 0.733833
R13793 nEN.n1139 nEN.n184 0.733833
R13794 nEN.n225 nEN.n222 0.573769
R13795 nEN.n281 nEN.n278 0.573769
R13796 nEN.n238 nEN.n235 0.573695
R13797 nEN.n292 nEN.n290 0.573695
R13798 nEN.n250 nEN.n247 0.573346
R13799 nEN.n1015 nEN.n236 0.573297
R13800 nEN.n717 nEN.n379 0.550549
R13801 nEN.n317 nEN.n316 0.550549
R13802 nEN.n1062 nEN.n221 0.39244
R13803 nEN.n954 nEN.n277 0.39244
R13804 nEN.n1037 nEN.n234 0.389994
R13805 nEN.n929 nEN.n291 0.389994
R13806 nEN.n1011 nEN.n246 0.387191
R13807 nEN.n1089 nEN.n206 0.384705
R13808 nEN.n989 nEN.n988 0.384705
R13809 nEN.n1064 nEN.n1063 0.384705
R13810 nEN.n955 nEN.n274 0.384705
R13811 nEN.n1088 nEN.n209 0.382331
R13812 nEN.n986 nEN.n260 0.382331
R13813 nEN.n1070 nEN.n210 0.382034
R13814 nEN.n962 nEN.n261 0.382034
R13815 nEN.n1044 nEN.n223 0.379547
R13816 nEN.n1002 nEN.n248 0.379547
R13817 nEN.n938 nEN.n279 0.379547
R13818 nEN.n1042 nEN.n223 0.375976
R13819 nEN.n940 nEN.n279 0.375976
R13820 nEN.n252 nEN.n248 0.375884
R13821 nEN.n1068 nEN.n210 0.374982
R13822 nEN.n964 nEN.n261 0.374982
R13823 nEN.n1088 nEN.n207 0.374889
R13824 nEN.n986 nEN.n259 0.374889
R13825 nEN.n1096 nEN.n1089 0.373984
R13826 nEN.n988 nEN.n256 0.373984
R13827 nEN.n1063 nEN.n220 0.373891
R13828 nEN.n956 nEN.n955 0.373891
R13829 nEN.n1019 nEN.n236 0.280767
R13830 nEN.n1127 nEN.n184 0.275034
R13831 nEN nEN.n1374 0.115637
R13832 nEN.n1375 nEN 0.106395
R13833 nEN.n917 nEN.n299 0.0405
R13834 nEN.n895 nEN.n299 0.0405
R13835 nEN.n895 nEN.n335 0.0405
R13836 nEN.n891 nEN.n335 0.0405
R13837 nEN.n891 nEN.n890 0.0405
R13838 nEN.n890 nEN.n889 0.0405
R13839 nEN.n889 nEN.n340 0.0405
R13840 nEN.n885 nEN.n340 0.0405
R13841 nEN.n885 nEN.n884 0.0405
R13842 nEN.n884 nEN.n883 0.0405
R13843 nEN.n883 nEN.n345 0.0405
R13844 nEN.n879 nEN.n345 0.0405
R13845 nEN.n879 nEN.n878 0.0405
R13846 nEN.n878 nEN.n877 0.0405
R13847 nEN.n873 nEN.n350 0.0405
R13848 nEN.n873 nEN.n872 0.0405
R13849 nEN.n872 nEN.n871 0.0405
R13850 nEN.n871 nEN.n355 0.0405
R13851 nEN.n867 nEN.n355 0.0405
R13852 nEN.n867 nEN.n866 0.0405
R13853 nEN.n866 nEN.n865 0.0405
R13854 nEN.n865 nEN.n360 0.0405
R13855 nEN.n861 nEN.n360 0.0405
R13856 nEN.n861 nEN.n860 0.0405
R13857 nEN.n860 nEN.n859 0.0405
R13858 nEN.n859 nEN.n365 0.0405
R13859 nEN.n1153 nEN.n168 0.0405
R13860 nEN.n1154 nEN.n1153 0.0405
R13861 nEN.n1155 nEN.n1154 0.0405
R13862 nEN.n1155 nEN.n156 0.0405
R13863 nEN.n1173 nEN.n156 0.0405
R13864 nEN.n1174 nEN.n1173 0.0405
R13865 nEN.n1175 nEN.n1174 0.0405
R13866 nEN.n1175 nEN.n143 0.0405
R13867 nEN.n1198 nEN.n143 0.0405
R13868 nEN.n1199 nEN.n1198 0.0405
R13869 nEN.n1200 nEN.n1199 0.0405
R13870 nEN.n1200 nEN.n132 0.0405
R13871 nEN.n1226 nEN.n132 0.0405
R13872 nEN.n1227 nEN.n1226 0.0405
R13873 nEN.n1228 nEN.n120 0.0405
R13874 nEN.n1246 nEN.n120 0.0405
R13875 nEN.n1247 nEN.n1246 0.0405
R13876 nEN.n1248 nEN.n1247 0.0405
R13877 nEN.n1248 nEN.n109 0.0405
R13878 nEN.n1275 nEN.n109 0.0405
R13879 nEN.n1276 nEN.n1275 0.0405
R13880 nEN.n1277 nEN.n1276 0.0405
R13881 nEN.n1277 nEN.n100 0.0405
R13882 nEN.n1299 nEN.n100 0.0405
R13883 nEN.n1300 nEN.n1299 0.0405
R13884 nEN.n1302 nEN.n1300 0.0405
R13885 nEN.n1152 nEN.n169 0.0405
R13886 nEN.n1152 nEN.n167 0.0405
R13887 nEN.n1156 nEN.n167 0.0405
R13888 nEN.n1156 nEN.n157 0.0405
R13889 nEN.n1172 nEN.n157 0.0405
R13890 nEN.n1172 nEN.n155 0.0405
R13891 nEN.n1176 nEN.n155 0.0405
R13892 nEN.n1176 nEN.n144 0.0405
R13893 nEN.n1197 nEN.n144 0.0405
R13894 nEN.n1197 nEN.n142 0.0405
R13895 nEN.n1201 nEN.n142 0.0405
R13896 nEN.n1201 nEN.n133 0.0405
R13897 nEN.n1225 nEN.n133 0.0405
R13898 nEN.n1225 nEN.n131 0.0405
R13899 nEN.n1229 nEN.n121 0.0405
R13900 nEN.n1245 nEN.n121 0.0405
R13901 nEN.n1245 nEN.n119 0.0405
R13902 nEN.n1249 nEN.n119 0.0405
R13903 nEN.n1249 nEN.n110 0.0405
R13904 nEN.n1274 nEN.n110 0.0405
R13905 nEN.n1274 nEN.n108 0.0405
R13906 nEN.n1278 nEN.n108 0.0405
R13907 nEN.n1278 nEN.n101 0.0405
R13908 nEN.n1298 nEN.n101 0.0405
R13909 nEN.n1298 nEN.n99 0.0405
R13910 nEN.n1303 nEN.n99 0.0405
R13911 nEN.n918 nEN.n298 0.0405
R13912 nEN.n894 nEN.n298 0.0405
R13913 nEN.n894 nEN.n893 0.0405
R13914 nEN.n893 nEN.n892 0.0405
R13915 nEN.n892 nEN.n336 0.0405
R13916 nEN.n888 nEN.n336 0.0405
R13917 nEN.n888 nEN.n887 0.0405
R13918 nEN.n887 nEN.n886 0.0405
R13919 nEN.n886 nEN.n341 0.0405
R13920 nEN.n882 nEN.n341 0.0405
R13921 nEN.n882 nEN.n881 0.0405
R13922 nEN.n881 nEN.n880 0.0405
R13923 nEN.n880 nEN.n346 0.0405
R13924 nEN.n876 nEN.n346 0.0405
R13925 nEN.n875 nEN.n874 0.0405
R13926 nEN.n874 nEN.n351 0.0405
R13927 nEN.n870 nEN.n351 0.0405
R13928 nEN.n870 nEN.n869 0.0405
R13929 nEN.n869 nEN.n868 0.0405
R13930 nEN.n868 nEN.n356 0.0405
R13931 nEN.n864 nEN.n356 0.0405
R13932 nEN.n864 nEN.n863 0.0405
R13933 nEN.n863 nEN.n862 0.0405
R13934 nEN.n862 nEN.n361 0.0405
R13935 nEN.n858 nEN.n361 0.0405
R13936 nEN.n858 nEN.n857 0.0405
R13937 nEN.n877 nEN.n350 0.0360676
R13938 nEN.n19 nEN.n3 0.0360676
R13939 nEN.n20 nEN.n19 0.0360676
R13940 nEN.n21 nEN.n20 0.0360676
R13941 nEN.n34 nEN.n21 0.0360676
R13942 nEN.n36 nEN.n34 0.0360676
R13943 nEN.n37 nEN.n36 0.0360676
R13944 nEN.n38 nEN.n37 0.0360676
R13945 nEN.n39 nEN.n38 0.0360676
R13946 nEN.n63 nEN.n39 0.0360676
R13947 nEN.n64 nEN.n63 0.0360676
R13948 nEN.n65 nEN.n64 0.0360676
R13949 nEN.n66 nEN.n65 0.0360676
R13950 nEN.n83 nEN.n66 0.0360676
R13951 nEN.n84 nEN.n83 0.0360676
R13952 nEN.n85 nEN.n84 0.0360676
R13953 nEN.n86 nEN.n85 0.0360676
R13954 nEN.n1228 nEN.n1227 0.0360676
R13955 nEN.n1229 nEN.n131 0.0360676
R13956 nEN.n922 nEN.n297 0.0360676
R13957 nEN.n297 nEN.n285 0.0360676
R13958 nEN.n944 nEN.n285 0.0360676
R13959 nEN.n944 nEN.n283 0.0360676
R13960 nEN.n948 nEN.n283 0.0360676
R13961 nEN.n948 nEN.n271 0.0360676
R13962 nEN.n968 nEN.n271 0.0360676
R13963 nEN.n968 nEN.n268 0.0360676
R13964 nEN.n979 nEN.n268 0.0360676
R13965 nEN.n979 nEN.n269 0.0360676
R13966 nEN.n975 nEN.n269 0.0360676
R13967 nEN.n975 nEN.n974 0.0360676
R13968 nEN.n974 nEN.n973 0.0360676
R13969 nEN.n973 nEN.n242 0.0360676
R13970 nEN.n1024 nEN.n242 0.0360676
R13971 nEN.n1024 nEN.n240 0.0360676
R13972 nEN.n1028 nEN.n240 0.0360676
R13973 nEN.n1028 nEN.n229 0.0360676
R13974 nEN.n1048 nEN.n229 0.0360676
R13975 nEN.n1048 nEN.n227 0.0360676
R13976 nEN.n1052 nEN.n227 0.0360676
R13977 nEN.n1052 nEN.n216 0.0360676
R13978 nEN.n1074 nEN.n216 0.0360676
R13979 nEN.n1074 nEN.n214 0.0360676
R13980 nEN.n1078 nEN.n214 0.0360676
R13981 nEN.n1078 nEN.n203 0.0360676
R13982 nEN.n1100 nEN.n203 0.0360676
R13983 nEN.n1100 nEN.n200 0.0360676
R13984 nEN.n1105 nEN.n200 0.0360676
R13985 nEN.n1105 nEN.n201 0.0360676
R13986 nEN.n201 nEN.n187 0.0360676
R13987 nEN.n1134 nEN.n187 0.0360676
R13988 nEN.n1134 nEN.n185 0.0360676
R13989 nEN.n921 nEN.n920 0.0360676
R13990 nEN.n920 nEN.n284 0.0360676
R13991 nEN.n945 nEN.n284 0.0360676
R13992 nEN.n946 nEN.n945 0.0360676
R13993 nEN.n947 nEN.n946 0.0360676
R13994 nEN.n947 nEN.n270 0.0360676
R13995 nEN.n969 nEN.n270 0.0360676
R13996 nEN.n970 nEN.n969 0.0360676
R13997 nEN.n978 nEN.n970 0.0360676
R13998 nEN.n978 nEN.n977 0.0360676
R13999 nEN.n977 nEN.n976 0.0360676
R14000 nEN.n976 nEN.n971 0.0360676
R14001 nEN.n972 nEN.n971 0.0360676
R14002 nEN.n972 nEN.n241 0.0360676
R14003 nEN.n1025 nEN.n241 0.0360676
R14004 nEN.n1026 nEN.n1025 0.0360676
R14005 nEN.n1027 nEN.n1026 0.0360676
R14006 nEN.n1027 nEN.n228 0.0360676
R14007 nEN.n1049 nEN.n228 0.0360676
R14008 nEN.n1050 nEN.n1049 0.0360676
R14009 nEN.n1051 nEN.n1050 0.0360676
R14010 nEN.n1051 nEN.n215 0.0360676
R14011 nEN.n1075 nEN.n215 0.0360676
R14012 nEN.n1076 nEN.n1075 0.0360676
R14013 nEN.n1077 nEN.n1076 0.0360676
R14014 nEN.n1077 nEN.n202 0.0360676
R14015 nEN.n1101 nEN.n202 0.0360676
R14016 nEN.n1102 nEN.n1101 0.0360676
R14017 nEN.n1104 nEN.n1102 0.0360676
R14018 nEN.n1104 nEN.n1103 0.0360676
R14019 nEN.n1103 nEN.n186 0.0360676
R14020 nEN.n1135 nEN.n186 0.0360676
R14021 nEN.n1136 nEN.n1135 0.0360676
R14022 nEN.n876 nEN.n875 0.0360676
R14023 nEN.n729 nEN.n366 0.0360676
R14024 nEN.n730 nEN.n729 0.0360676
R14025 nEN.n731 nEN.n730 0.0360676
R14026 nEN.n744 nEN.n731 0.0360676
R14027 nEN.n746 nEN.n744 0.0360676
R14028 nEN.n747 nEN.n746 0.0360676
R14029 nEN.n748 nEN.n747 0.0360676
R14030 nEN.n749 nEN.n748 0.0360676
R14031 nEN.n773 nEN.n749 0.0360676
R14032 nEN.n774 nEN.n773 0.0360676
R14033 nEN.n775 nEN.n774 0.0360676
R14034 nEN.n776 nEN.n775 0.0360676
R14035 nEN.n777 nEN.n776 0.0360676
R14036 nEN.n777 nEN.n4 0.0360676
R14037 nEN.n854 nEN.n368 0.0360676
R14038 nEN.n842 nEN.n368 0.0360676
R14039 nEN.n842 nEN.n841 0.0360676
R14040 nEN.n841 nEN.n732 0.0360676
R14041 nEN.n745 nEN.n732 0.0360676
R14042 nEN.n745 nEN.n743 0.0360676
R14043 nEN.n825 nEN.n743 0.0360676
R14044 nEN.n825 nEN.n824 0.0360676
R14045 nEN.n824 nEN.n750 0.0360676
R14046 nEN.n772 nEN.n750 0.0360676
R14047 nEN.n812 nEN.n772 0.0360676
R14048 nEN.n812 nEN.n811 0.0360676
R14049 nEN.n811 nEN.n778 0.0360676
R14050 nEN.n791 nEN.n778 0.0360676
R14051 nEN.n791 nEN.n5 0.0360676
R14052 nEN.n1372 nEN.n1371 0.0360676
R14053 nEN.n1371 nEN.n7 0.0360676
R14054 nEN.n1360 nEN.n7 0.0360676
R14055 nEN.n1360 nEN.n1359 0.0360676
R14056 nEN.n1359 nEN.n22 0.0360676
R14057 nEN.n35 nEN.n22 0.0360676
R14058 nEN.n35 nEN.n33 0.0360676
R14059 nEN.n1343 nEN.n33 0.0360676
R14060 nEN.n1343 nEN.n1342 0.0360676
R14061 nEN.n1342 nEN.n40 0.0360676
R14062 nEN.n62 nEN.n40 0.0360676
R14063 nEN.n1330 nEN.n62 0.0360676
R14064 nEN.n1330 nEN.n1329 0.0360676
R14065 nEN.n1329 nEN.n67 0.0360676
R14066 nEN.n82 nEN.n67 0.0360676
R14067 nEN.n1317 nEN.n82 0.0360676
R14068 nEN.n1317 nEN.n1316 0.0360676
R14069 nEN.n917 nEN.n296 0.0234189
R14070 nEN.n1137 nEN.n168 0.0234189
R14071 nEN.n1138 nEN.n169 0.0234189
R14072 nEN.n919 nEN.n918 0.0234189
R14073 nEN.n855 nEN.n365 0.0233108
R14074 nEN.n1302 nEN.n1301 0.0233108
R14075 nEN.n1303 nEN.n87 0.0233108
R14076 nEN.n857 nEN.n856 0.0233108
R14077 nEN.n922 nEN.n296 0.0227703
R14078 nEN.n921 nEN.n919 0.0227703
R14079 nEN.n856 nEN.n366 0.0227703
R14080 nEN.n855 nEN.n854 0.0227703
R14081 nEN.n897 nEN.n330 0.0188784
R14082 nEN.n473 nEN.n334 0.0188784
R14083 nEN.n482 nEN.n481 0.0188784
R14084 nEN.n491 nEN.n490 0.0188784
R14085 nEN.n498 nEN.n497 0.0188784
R14086 nEN.n524 nEN.n523 0.0188784
R14087 nEN.n532 nEN.n531 0.0188784
R14088 nEN.n539 nEN.n538 0.0188784
R14089 nEN.n554 nEN.n440 0.0188784
R14090 nEN.n557 nEN.n556 0.0188784
R14091 nEN.n571 nEN.n433 0.0188784
R14092 nEN.n581 nEN.n580 0.0188784
R14093 nEN.n590 nEN.n589 0.0188784
R14094 nEN.n599 nEN.n598 0.0188784
R14095 nEN.n608 nEN.n607 0.0188784
R14096 nEN.n615 nEN.n614 0.0188784
R14097 nEN.n626 nEN.n624 0.0188784
R14098 nEN.n640 nEN.n409 0.0188784
R14099 nEN.n656 nEN.n655 0.0188784
R14100 nEN.n671 nEN.n397 0.0188784
R14101 nEN.n674 nEN.n673 0.0188784
R14102 nEN.n682 nEN.n681 0.0188784
R14103 nEN.n690 nEN.n390 0.0188784
R14104 nEN.n178 nEN.n171 0.0188784
R14105 nEN.n176 nEN.n166 0.0188784
R14106 nEN.n1161 nEN.n1158 0.0188784
R14107 nEN.n1159 nEN.n158 0.0188784
R14108 nEN.n1170 nEN.n160 0.0188784
R14109 nEN.n1184 nEN.n1183 0.0188784
R14110 nEN.n1186 nEN.n145 0.0188784
R14111 nEN.n1195 nEN.n147 0.0188784
R14112 nEN.n1203 nEN.n141 0.0188784
R14113 nEN.n1208 nEN.n139 0.0188784
R14114 nEN.n1211 nEN.n1210 0.0188784
R14115 nEN.n1223 nEN.n135 0.0188784
R14116 nEN.n1219 nEN.n130 0.0188784
R14117 nEN.n1234 nEN.n1231 0.0188784
R14118 nEN.n1232 nEN.n122 0.0188784
R14119 nEN.n1243 nEN.n124 0.0188784
R14120 nEN.n1251 nEN.n118 0.0188784
R14121 nEN.n1256 nEN.n116 0.0188784
R14122 nEN.n1272 nEN.n112 0.0188784
R14123 nEN.n1267 nEN.n107 0.0188784
R14124 nEN.n1283 nEN.n1280 0.0188784
R14125 nEN.n1281 nEN.n102 0.0188784
R14126 nEN.n1296 nEN.n103 0.0188784
R14127 nEN.n369 nEN.n367 0.0188784
R14128 nEN.n852 nEN.n370 0.0188784
R14129 nEN.n844 nEN.n727 0.0188784
R14130 nEN.n733 nEN.n728 0.0188784
R14131 nEN.n795 nEN.n8 0.0188784
R14132 nEN.n1369 nEN.n9 0.0188784
R14133 nEN.n1362 nEN.n17 0.0188784
R14134 nEN.n23 nEN.n18 0.0188784
R14135 nEN.n305 nEN.n295 0.0188784
R14136 nEN.n925 nEN.n924 0.0188784
R14137 nEN.n934 nEN.n933 0.0188784
R14138 nEN.n936 nEN.n286 0.0188784
R14139 nEN.n1017 nEN.n239 0.0188784
R14140 nEN.n1033 nEN.n1030 0.0188784
R14141 nEN.n1031 nEN.n230 0.0188784
R14142 nEN.n1046 nEN.n232 0.0188784
R14143 nEN.n915 nEN.n301 0.0187703
R14144 nEN.n330 nEN.n329 0.0187703
R14145 nEN.n509 nEN.n507 0.0187703
R14146 nEN.n523 nEN.n452 0.0187703
R14147 nEN.n572 nEN.n571 0.0187703
R14148 nEN.n641 nEN.n640 0.0187703
R14149 nEN.n649 nEN.n648 0.0187703
R14150 nEN.n390 nEN.n389 0.0187703
R14151 nEN.n709 nEN.n382 0.0187703
R14152 nEN.n1142 nEN.n170 0.0187703
R14153 nEN.n1150 nEN.n171 0.0187703
R14154 nEN.n1178 nEN.n154 0.0187703
R14155 nEN.n1183 nEN.n152 0.0187703
R14156 nEN.n1211 nEN.n134 0.0187703
R14157 nEN.n1257 nEN.n1256 0.0187703
R14158 nEN.n1259 nEN.n111 0.0187703
R14159 nEN.n1291 nEN.n103 0.0187703
R14160 nEN.n1305 nEN.n98 0.0187703
R14161 nEN.n836 nEN.n835 0.0187703
R14162 nEN.n832 nEN.n831 0.0187703
R14163 nEN.n828 nEN.n827 0.0187703
R14164 nEN.n751 nEN.n742 0.0187703
R14165 nEN.n822 nEN.n752 0.0187703
R14166 nEN.n770 nEN.n768 0.0187703
R14167 nEN.n814 nEN.n765 0.0187703
R14168 nEN.n779 nEN.n766 0.0187703
R14169 nEN.n809 nEN.n780 0.0187703
R14170 nEN.n790 nEN.n789 0.0187703
R14171 nEN.n802 nEN.n801 0.0187703
R14172 nEN.n799 nEN.n793 0.0187703
R14173 nEN.n1354 nEN.n1353 0.0187703
R14174 nEN.n1350 nEN.n1349 0.0187703
R14175 nEN.n1346 nEN.n1345 0.0187703
R14176 nEN.n41 nEN.n32 0.0187703
R14177 nEN.n1340 nEN.n42 0.0187703
R14178 nEN.n60 nEN.n58 0.0187703
R14179 nEN.n1332 nEN.n55 0.0187703
R14180 nEN.n68 nEN.n56 0.0187703
R14181 nEN.n1327 nEN.n69 0.0187703
R14182 nEN.n79 nEN.n78 0.0187703
R14183 nEN.n1320 nEN.n1319 0.0187703
R14184 nEN.n88 nEN.n81 0.0187703
R14185 nEN.n950 nEN.n282 0.0187703
R14186 nEN.n958 nEN.n275 0.0187703
R14187 nEN.n960 nEN.n272 0.0187703
R14188 nEN.n966 nEN.n273 0.0187703
R14189 nEN.n982 nEN.n981 0.0187703
R14190 nEN.n267 nEN.n265 0.0187703
R14191 nEN.n992 nEN.n991 0.0187703
R14192 nEN.n996 nEN.n995 0.0187703
R14193 nEN.n1000 nEN.n999 0.0187703
R14194 nEN.n1005 nEN.n1004 0.0187703
R14195 nEN.n1007 nEN.n243 0.0187703
R14196 nEN.n1022 nEN.n244 0.0187703
R14197 nEN.n1058 nEN.n1054 0.0187703
R14198 nEN.n1056 nEN.n217 0.0187703
R14199 nEN.n1072 nEN.n218 0.0187703
R14200 nEN.n1066 nEN.n213 0.0187703
R14201 nEN.n1084 nEN.n1083 0.0187703
R14202 nEN.n1081 nEN.n204 0.0187703
R14203 nEN.n1098 nEN.n205 0.0187703
R14204 nEN.n1093 nEN.n199 0.0187703
R14205 nEN.n1108 nEN.n1107 0.0187703
R14206 nEN.n1121 nEN.n1118 0.0187703
R14207 nEN.n1119 nEN.n188 0.0187703
R14208 nEN.n1132 nEN.n189 0.0187703
R14209 nEN.n1373 nEN.n1372 0.0186443
R14210 nEN.n1373 nEN.n5 0.0186443
R14211 nEN.n896 nEN.n334 0.0185541
R14212 nEN.n681 nEN.n363 0.0185541
R14213 nEN.n177 nEN.n176 0.0185541
R14214 nEN.n1297 nEN.n102 0.0185541
R14215 nEN.n839 nEN.n734 0.0184459
R14216 nEN.n1357 nEN.n24 0.0184459
R14217 nEN.n942 nEN.n287 0.0184459
R14218 nEN.n1053 nEN.n226 0.0184459
R14219 nEN.n580 nEN.n348 0.0182297
R14220 nEN.n1224 nEN.n1223 0.0182297
R14221 nEN.n840 nEN.n839 0.0181216
R14222 nEN.n1358 nEN.n1357 0.0181216
R14223 nEN.n943 nEN.n942 0.0181216
R14224 nEN.n231 nEN.n226 0.0181216
R14225 nEN.n509 nEN.n508 0.0175811
R14226 nEN.n648 nEN.n357 0.0175811
R14227 nEN.n1178 nEN.n1177 0.0175811
R14228 nEN.n1259 nEN.n1258 0.0175811
R14229 nEN.n835 nEN.n738 0.0173649
R14230 nEN.n1353 nEN.n28 0.0173649
R14231 nEN.n950 nEN.n949 0.0173649
R14232 nEN.n1058 nEN.n1057 0.0173649
R14233 nEN.n843 nEN.n728 0.0170405
R14234 nEN.n1361 nEN.n18 0.0170405
R14235 nEN.n936 nEN.n935 0.0170405
R14236 nEN.n1047 nEN.n1046 0.0170405
R14237 nEN.n531 nEN.n342 0.0167162
R14238 nEN.n626 nEN.n625 0.0167162
R14239 nEN.n1186 nEN.n1185 0.0167162
R14240 nEN.n1251 nEN.n1250 0.0167162
R14241 nEN.n831 nEN.n740 0.0162838
R14242 nEN.n1349 nEN.n30 0.0162838
R14243 nEN.n959 nEN.n958 0.0162838
R14244 nEN.n1073 nEN.n217 0.0162838
R14245 nEN.n556 nEN.n347 0.0159595
R14246 nEN.n598 nEN.n422 0.0159595
R14247 nEN.n1209 nEN.n1208 0.0159595
R14248 nEN.n1231 nEN.n1230 0.0159595
R14249 nEN.n727 nEN.n726 0.0159595
R14250 nEN.n17 nEN.n16 0.0159595
R14251 nEN.n933 nEN.n289 0.0159595
R14252 nEN.n1032 nEN.n1031 0.0159595
R14253 nEN.n328 nEN.n301 0.0157432
R14254 nEN.n382 nEN.n364 0.0157432
R14255 nEN.n1151 nEN.n170 0.0157432
R14256 nEN.n1290 nEN.n98 0.0157432
R14257 nEN.n481 nEN.n465 0.0152027
R14258 nEN.n673 nEN.n362 0.0152027
R14259 nEN.n1158 nEN.n1157 0.0152027
R14260 nEN.n1283 nEN.n1282 0.0152027
R14261 nEN.n827 nEN.n826 0.0152027
R14262 nEN.n1345 nEN.n1344 0.0152027
R14263 nEN.n967 nEN.n272 0.0152027
R14264 nEN.n1065 nEN.n218 0.0152027
R14265 nEN.n589 nEN.n349 0.0148784
R14266 nEN.n1219 nEN.n1218 0.0148784
R14267 nEN.n853 nEN.n852 0.0148784
R14268 nEN.n1370 nEN.n1369 0.0148784
R14269 nEN.n924 nEN.n923 0.0148784
R14270 nEN.n1030 nEN.n1029 0.0148784
R14271 nEN.n497 nEN.n339 0.0141216
R14272 nEN.n655 nEN.n358 0.0141216
R14273 nEN.n160 nEN.n159 0.0141216
R14274 nEN.n1273 nEN.n1272 0.0141216
R14275 nEN.n823 nEN.n751 0.0141216
R14276 nEN.n1341 nEN.n41 0.0141216
R14277 nEN.n273 nEN.n264 0.0141216
R14278 nEN.n1079 nEN.n213 0.0141216
R14279 nEN.n1301 nEN.n86 0.0137973
R14280 nEN.n795 nEN.n6 0.0137973
R14281 nEN.n1315 nEN.n1314 0.0137973
R14282 nEN.n1017 nEN.n1016 0.0137973
R14283 nEN.n1139 nEN.n182 0.0137973
R14284 nEN.n1138 nEN.n185 0.0137973
R14285 nEN.n1137 nEN.n1136 0.0137973
R14286 nEN.n1316 nEN.n87 0.0137973
R14287 nEN.n1312 nEN.n73 0.0134381
R14288 nEN.n538 nEN.n343 0.0133649
R14289 nEN.n614 nEN.n354 0.0133649
R14290 nEN.n1196 nEN.n1195 0.0133649
R14291 nEN.n124 nEN.n123 0.0133649
R14292 nEN.n767 nEN.n752 0.0130405
R14293 nEN.n57 nEN.n42 0.0130405
R14294 nEN.n981 nEN.n980 0.0130405
R14295 nEN.n1083 nEN.n1082 0.0130405
R14296 nEN.n800 nEN.n799 0.0128243
R14297 nEN.n1318 nEN.n81 0.0128243
R14298 nEN.n1023 nEN.n1022 0.0128243
R14299 nEN.n1133 nEN.n1132 0.0128243
R14300 nEN.n555 nEN.n554 0.0126081
R14301 nEN.n607 nEN.n352 0.0126081
R14302 nEN.n1203 nEN.n1202 0.0126081
R14303 nEN.n1233 nEN.n1232 0.0126081
R14304 nEN.n916 nEN.n300 0.0123919
R14305 nEN.n711 nEN.n710 0.0123919
R14306 nEN.n1141 nEN.n1140 0.0123919
R14307 nEN.n1304 nEN.n89 0.0123919
R14308 nEN.n771 nEN.n770 0.0119595
R14309 nEN.n61 nEN.n60 0.0119595
R14310 nEN.n265 nEN.n257 0.0119595
R14311 nEN.n1099 nEN.n204 0.0119595
R14312 nEN.n490 nEN.n337 0.0118514
R14313 nEN.n672 nEN.n671 0.0118514
R14314 nEN.n1160 nEN.n1159 0.0118514
R14315 nEN.n1279 nEN.n107 0.0118514
R14316 nEN.n802 nEN.n792 0.0117432
R14317 nEN.n1320 nEN.n80 0.0117432
R14318 nEN.n1007 nEN.n1006 0.0117432
R14319 nEN.n1120 nEN.n1119 0.0117432
R14320 nEN.n1127 nEN.n180 0.0116588
R14321 nEN.n305 nEN.n300 0.011527
R14322 nEN.n1140 nEN.n1139 0.011527
R14323 nEN.n711 nEN.n367 0.0114189
R14324 nEN.n1314 nEN.n89 0.0114189
R14325 nEN.n930 nEN.n279 0.0109762
R14326 nEN.n955 nEN.n954 0.0109762
R14327 nEN.n985 nEN.n261 0.0109762
R14328 nEN.n988 nEN.n986 0.0109762
R14329 nEN.n987 nEN.n248 0.0109762
R14330 nEN.n1012 nEN.n1011 0.0109762
R14331 nEN.n1037 nEN.n236 0.0109762
R14332 nEN.n1038 nEN.n223 0.0109762
R14333 nEN.n1063 nEN.n1062 0.0109762
R14334 nEN.n1087 nEN.n210 0.0109762
R14335 nEN.n1089 nEN.n1088 0.0109762
R14336 nEN.n1146 nEN.n1145 0.0109762
R14337 nEN.n1146 nEN.n162 0.0109762
R14338 nEN.n1164 nEN.n162 0.0109762
R14339 nEN.n1165 nEN.n1164 0.0109762
R14340 nEN.n1166 nEN.n1165 0.0109762
R14341 nEN.n1166 nEN.n149 0.0109762
R14342 nEN.n1189 nEN.n149 0.0109762
R14343 nEN.n1190 nEN.n1189 0.0109762
R14344 nEN.n1191 nEN.n1190 0.0109762
R14345 nEN.n1191 nEN.n137 0.0109762
R14346 nEN.n1214 nEN.n137 0.0109762
R14347 nEN.n1215 nEN.n126 0.0109762
R14348 nEN.n1237 nEN.n126 0.0109762
R14349 nEN.n1238 nEN.n1237 0.0109762
R14350 nEN.n1239 nEN.n1238 0.0109762
R14351 nEN.n1239 nEN.n114 0.0109762
R14352 nEN.n1262 nEN.n114 0.0109762
R14353 nEN.n1263 nEN.n1262 0.0109762
R14354 nEN.n1263 nEN.n105 0.0109762
R14355 nEN.n1286 nEN.n105 0.0109762
R14356 nEN.n1287 nEN.n1286 0.0109762
R14357 nEN.n1287 nEN.n96 0.0109762
R14358 nEN.n1308 nEN.n96 0.0109762
R14359 nEN.n847 nEN.n723 0.0109762
R14360 nEN.n756 nEN.n755 0.0109762
R14361 nEN.n761 nEN.n760 0.0109762
R14362 nEN.n818 nEN.n817 0.0109762
R14363 nEN.n806 nEN.n762 0.0109762
R14364 nEN.n805 nEN.n784 0.0109762
R14365 nEN.n1366 nEN.n12 0.0109762
R14366 nEN.n1365 nEN.n13 0.0109762
R14367 nEN.n46 nEN.n45 0.0109762
R14368 nEN.n51 nEN.n50 0.0109762
R14369 nEN.n1336 nEN.n1335 0.0109762
R14370 nEN.n1324 nEN.n52 0.0109762
R14371 nEN.n1323 nEN.n73 0.0109762
R14372 nEN.n930 nEN.n929 0.01095
R14373 nEN.n954 nEN.n279 0.01095
R14374 nEN.n955 nEN.n261 0.01095
R14375 nEN.n986 nEN.n985 0.01095
R14376 nEN.n988 nEN.n987 0.01095
R14377 nEN.n1011 nEN.n248 0.01095
R14378 nEN.n1012 nEN.n236 0.01095
R14379 nEN.n1038 nEN.n1037 0.01095
R14380 nEN.n1062 nEN.n223 0.01095
R14381 nEN.n1063 nEN.n210 0.01095
R14382 nEN.n1088 nEN.n1087 0.01095
R14383 nEN.n1090 nEN.n1089 0.01095
R14384 nEN.n1215 nEN.n1214 0.01095
R14385 nEN.n1309 nEN.n1308 0.01095
R14386 nEN.n755 nEN.n723 0.01095
R14387 nEN.n760 nEN.n756 0.01095
R14388 nEN.n818 nEN.n761 0.01095
R14389 nEN.n817 nEN.n762 0.01095
R14390 nEN.n806 nEN.n805 0.01095
R14391 nEN.n784 nEN.n12 0.01095
R14392 nEN.n1366 nEN.n1365 0.01095
R14393 nEN.n45 nEN.n13 0.01095
R14394 nEN.n50 nEN.n46 0.01095
R14395 nEN.n1336 nEN.n51 0.01095
R14396 nEN.n1335 nEN.n52 0.01095
R14397 nEN.n1324 nEN.n1323 0.01095
R14398 nEN.n814 nEN.n813 0.0108784
R14399 nEN.n1332 nEN.n1331 0.0108784
R14400 nEN.n992 nEN.n255 0.0108784
R14401 nEN.n1092 nEN.n205 0.0108784
R14402 nEN.n491 nEN.n338 0.0107703
R14403 nEN.n397 nEN.n359 0.0107703
R14404 nEN.n1171 nEN.n158 0.0107703
R14405 nEN.n1267 nEN.n1266 0.0107703
R14406 nEN.n789 nEN.n787 0.0106622
R14407 nEN.n78 nEN.n76 0.0106622
R14408 nEN.n1004 nEN.n251 0.0106622
R14409 nEN.n1118 nEN.n195 0.0106622
R14410 nEN.n1145 nEN.n180 0.0106095
R14411 nEN.n440 nEN.n344 0.0100135
R14412 nEN.n608 nEN.n353 0.0100135
R14413 nEN.n146 nEN.n141 0.0100135
R14414 nEN.n1244 nEN.n122 0.0100135
R14415 nEN.n810 nEN.n779 0.0097973
R14416 nEN.n1328 nEN.n68 0.0097973
R14417 nEN.n996 nEN.n253 0.0097973
R14418 nEN.n1106 nEN.n199 0.0097973
R14419 nEN.n1128 nEN.n1127 0.00967266
R14420 nEN.n810 nEN.n809 0.00958108
R14421 nEN.n1328 nEN.n1327 0.00958108
R14422 nEN.n999 nEN.n253 0.00958108
R14423 nEN.n1108 nEN.n1106 0.00958108
R14424 nEN.n539 nEN.n344 0.00925676
R14425 nEN.n615 nEN.n353 0.00925676
R14426 nEN.n147 nEN.n146 0.00925676
R14427 nEN.n1244 nEN.n1243 0.00925676
R14428 nEN.n1011 nEN.n247 0.00880612
R14429 nEN.n787 nEN.n780 0.00871622
R14430 nEN.n76 nEN.n69 0.00871622
R14431 nEN.n1000 nEN.n251 0.00871622
R14432 nEN.n1107 nEN.n195 0.00871622
R14433 nEN.n498 nEN.n338 0.0085
R14434 nEN.n656 nEN.n359 0.0085
R14435 nEN.n1171 nEN.n1170 0.0085
R14436 nEN.n1266 nEN.n112 0.0085
R14437 nEN.n813 nEN.n766 0.0085
R14438 nEN.n1331 nEN.n56 0.0085
R14439 nEN.n995 nEN.n255 0.0085
R14440 nEN.n1093 nEN.n1092 0.0085
R14441 nEN.n1374 nEN.n3 0.00839189
R14442 nEN.n848 nEN.n847 0.00809524
R14443 nEN.n1126 nEN.n1125 0.00778095
R14444 nEN.n792 nEN.n790 0.00763514
R14445 nEN.n80 nEN.n79 0.00763514
R14446 nEN.n1006 nEN.n1005 0.00763514
R14447 nEN.n1121 nEN.n1120 0.00763514
R14448 nEN.n482 nEN.n337 0.00741892
R14449 nEN.n674 nEN.n672 0.00741892
R14450 nEN.n1161 nEN.n1160 0.00741892
R14451 nEN.n1280 nEN.n1279 0.00741892
R14452 nEN.n771 nEN.n765 0.00741892
R14453 nEN.n61 nEN.n55 0.00741892
R14454 nEN.n991 nEN.n257 0.00741892
R14455 nEN.n1099 nEN.n1098 0.00741892
R14456 nEN.n1090 nEN.n197 0.00725714
R14457 nEN.n1128 nEN.n1126 0.00707381
R14458 nEN.n916 nEN.n915 0.00698649
R14459 nEN.n710 nEN.n709 0.00698649
R14460 nEN.n1142 nEN.n1141 0.00698649
R14461 nEN.n1305 nEN.n1304 0.00698649
R14462 nEN.n929 nEN.n293 0.00696162
R14463 nEN.n1309 nEN.n95 0.00691667
R14464 nEN.n557 nEN.n555 0.00666216
R14465 nEN.n599 nEN.n352 0.00666216
R14466 nEN.n1202 nEN.n139 0.00666216
R14467 nEN.n1234 nEN.n1233 0.00666216
R14468 nEN.n801 nEN.n800 0.00655405
R14469 nEN.n1319 nEN.n1318 0.00655405
R14470 nEN.n1023 nEN.n243 0.00655405
R14471 nEN.n1133 nEN.n188 0.00655405
R14472 nEN.n768 nEN.n767 0.00633784
R14473 nEN.n58 nEN.n57 0.00633784
R14474 nEN.n980 nEN.n267 0.00633784
R14475 nEN.n1082 nEN.n1081 0.00633784
R14476 nEN.n532 nEN.n343 0.00590541
R14477 nEN.n624 nEN.n354 0.00590541
R14478 nEN.n1196 nEN.n145 0.00590541
R14479 nEN.n123 nEN.n118 0.00590541
R14480 nEN.n1037 nEN.n235 0.00588776
R14481 nEN.n929 nEN.n292 0.00588776
R14482 nEN.n793 nEN.n6 0.00547297
R14483 nEN.n1315 nEN.n88 0.00547297
R14484 nEN.n1016 nEN.n244 0.00547297
R14485 nEN.n189 nEN.n182 0.00547297
R14486 nEN.n823 nEN.n822 0.00525676
R14487 nEN.n1341 nEN.n1340 0.00525676
R14488 nEN.n982 nEN.n264 0.00525676
R14489 nEN.n1084 nEN.n1079 0.00525676
R14490 nEN.n507 nEN.n339 0.00514865
R14491 nEN.n649 nEN.n358 0.00514865
R14492 nEN.n159 nEN.n154 0.00514865
R14493 nEN.n1273 nEN.n111 0.00514865
R14494 nEN.n1312 nEN.n1311 0.00440238
R14495 nEN.n581 nEN.n349 0.00439189
R14496 nEN.n1218 nEN.n135 0.00439189
R14497 nEN.n853 nEN.n369 0.00439189
R14498 nEN.n1370 nEN.n8 0.00439189
R14499 nEN.n923 nEN.n295 0.00439189
R14500 nEN.n1029 nEN.n239 0.00439189
R14501 nEN.n1143 nEN.n181 0.00425921
R14502 nEN.n1149 nEN.n172 0.00425921
R14503 nEN.n165 nEN.n164 0.00425921
R14504 nEN.n1169 nEN.n1168 0.00425921
R14505 nEN.n1182 nEN.n150 0.00425921
R14506 nEN.n1187 nEN.n151 0.00425921
R14507 nEN.n1194 nEN.n1193 0.00425921
R14508 nEN.n1204 nEN.n140 0.00425921
R14509 nEN.n1222 nEN.n1221 0.00425921
R14510 nEN.n129 nEN.n128 0.00425921
R14511 nEN.n1242 nEN.n1241 0.00425921
R14512 nEN.n1252 nEN.n117 0.00425921
R14513 nEN.n1255 nEN.n1254 0.00425921
R14514 nEN.n1271 nEN.n1270 0.00425921
R14515 nEN.n1268 nEN.n1265 0.00425921
R14516 nEN.n1292 nEN.n97 0.00425921
R14517 nEN.n1306 nEN.n90 0.00425921
R14518 nEN.n735 nEN.n725 0.00425921
R14519 nEN.n838 nEN.n837 0.00425921
R14520 nEN.n834 nEN.n833 0.00425921
R14521 nEN.n830 nEN.n829 0.00425921
R14522 nEN.n769 nEN.n763 0.00425921
R14523 nEN.n815 nEN.n764 0.00425921
R14524 nEN.n808 nEN.n782 0.00425921
R14525 nEN.n788 nEN.n783 0.00425921
R14526 nEN.n796 nEN.n10 0.00425921
R14527 nEN.n25 nEN.n15 0.00425921
R14528 nEN.n1356 nEN.n1355 0.00425921
R14529 nEN.n1352 nEN.n1351 0.00425921
R14530 nEN.n1348 nEN.n1347 0.00425921
R14531 nEN.n59 nEN.n53 0.00425921
R14532 nEN.n1333 nEN.n54 0.00425921
R14533 nEN.n1326 nEN.n71 0.00425921
R14534 nEN.n77 nEN.n72 0.00425921
R14535 nEN.n994 nEN.n993 0.00425921
R14536 nEN.n998 nEN.n997 0.00425921
R14537 nEN.n1095 nEN.n1094 0.00425921
R14538 nEN.n1109 nEN.n198 0.00425921
R14539 nEN.n1115 nEN.n1113 0.00424524
R14540 nEN.n1149 nEN.n1148 0.0042371
R14541 nEN.n179 nEN.n175 0.0042371
R14542 nEN.n173 nEN.n163 0.0042371
R14543 nEN.n1162 nEN.n165 0.0042371
R14544 nEN.n1179 nEN.n153 0.0042371
R14545 nEN.n1182 nEN.n1181 0.0042371
R14546 nEN.n1205 nEN.n1204 0.0042371
R14547 nEN.n1207 nEN.n138 0.0042371
R14548 nEN.n1212 nEN.n136 0.0042371
R14549 nEN.n1222 nEN.n136 0.0042371
R14550 nEN.n1221 nEN.n1220 0.0042371
R14551 nEN.n1216 nEN.n127 0.0042371
R14552 nEN.n1235 nEN.n129 0.0042371
R14553 nEN.n1255 nEN.n115 0.0042371
R14554 nEN.n1260 nEN.n113 0.0042371
R14555 nEN.n1265 nEN.n106 0.0042371
R14556 nEN.n1284 nEN.n104 0.0042371
R14557 nEN.n1295 nEN.n1289 0.0042371
R14558 nEN.n1293 nEN.n1292 0.0042371
R14559 nEN.n724 nEN.n722 0.0042371
R14560 nEN.n845 nEN.n725 0.0042371
R14561 nEN.n829 nEN.n741 0.0042371
R14562 nEN.n758 nEN.n757 0.0042371
R14563 nEN.n821 nEN.n820 0.0042371
R14564 nEN.n769 nEN.n754 0.0042371
R14565 nEN.n788 nEN.n785 0.0042371
R14566 nEN.n803 nEN.n786 0.0042371
R14567 nEN.n798 nEN.n797 0.0042371
R14568 nEN.n797 nEN.n796 0.0042371
R14569 nEN.n1368 nEN.n10 0.0042371
R14570 nEN.n14 nEN.n11 0.0042371
R14571 nEN.n1363 nEN.n15 0.0042371
R14572 nEN.n1347 nEN.n31 0.0042371
R14573 nEN.n48 nEN.n47 0.0042371
R14574 nEN.n1339 nEN.n1338 0.0042371
R14575 nEN.n59 nEN.n44 0.0042371
R14576 nEN.n77 nEN.n74 0.0042371
R14577 nEN.n1321 nEN.n75 0.0042371
R14578 nEN.n93 nEN.n92 0.0042371
R14579 nEN.n1313 nEN.n93 0.0042371
R14580 nEN.n937 nEN.n288 0.0042371
R14581 nEN.n965 nEN.n262 0.0042371
R14582 nEN.n983 nEN.n263 0.0042371
R14583 nEN.n1021 nEN.n1020 0.0042371
R14584 nEN.n1045 nEN.n1040 0.0042371
R14585 nEN.n1067 nEN.n211 0.0042371
R14586 nEN.n1085 nEN.n212 0.0042371
R14587 nEN.n192 nEN.n191 0.0042371
R14588 nEN.n1131 nEN.n1130 0.0042371
R14589 nEN.n720 nEN.n719 0.00423273
R14590 nEN.n1020 nEN.n1019 0.00423268
R14591 nEN.n378 nEN.n375 0.00422178
R14592 nEN.n315 nEN.n314 0.00422178
R14593 nEN.n1112 nEN.n197 0.00421905
R14594 nEN.n826 nEN.n742 0.00417568
R14595 nEN.n1344 nEN.n32 0.00417568
R14596 nEN.n967 nEN.n966 0.00417568
R14597 nEN.n1066 nEN.n1065 0.00417568
R14598 nEN.n1147 nEN.n179 0.00410442
R14599 nEN.n1295 nEN.n1294 0.00410442
R14600 nEN.n473 nEN.n465 0.00406757
R14601 nEN.n682 nEN.n362 0.00406757
R14602 nEN.n1157 nEN.n166 0.00406757
R14603 nEN.n1282 nEN.n1281 0.00406757
R14604 nEN.n250 nEN.n245 0.00402269
R14605 nEN.n941 nEN.n277 0.00398793
R14606 nEN.n1041 nEN.n221 0.00398793
R14607 nEN.n838 nEN.n736 0.00397174
R14608 nEN.n808 nEN.n807 0.00397174
R14609 nEN.n1356 nEN.n26 0.00397174
R14610 nEN.n1326 nEN.n1325 0.00397174
R14611 nEN.n1193 nEN.n1192 0.00394963
R14612 nEN.n1242 nEN.n125 0.00394963
R14613 nEN.n932 nEN.n290 0.00394626
R14614 nEN.n238 nEN.n233 0.00394626
R14615 nEN.n309 nEN.n291 0.00393696
R14616 nEN.n1014 nEN.n234 0.00393696
R14617 nEN.n281 nEN.n276 0.00390294
R14618 nEN.n1055 nEN.n225 0.00390294
R14619 nEN.n1003 nEN.n246 0.00389381
R14620 nEN.n961 nEN.n274 0.00385851
R14621 nEN.n989 nEN.n258 0.00385851
R14622 nEN.n1071 nEN.n1064 0.00385851
R14623 nEN.n208 nEN.n206 0.00385851
R14624 nEN.n962 nEN.n961 0.00380768
R14625 nEN.n1071 nEN.n1070 0.00380768
R14626 nEN.n260 nEN.n258 0.00380053
R14627 nEN.n209 nEN.n208 0.00380053
R14628 nEN.n1169 nEN.n161 0.00379484
R14629 nEN.n1270 nEN.n1269 0.00379484
R14630 nEN.n718 nEN.n374 0.00379484
R14631 nEN.n1129 nEN.n184 0.00377273
R14632 nEN.n938 nEN.n937 0.0037725
R14633 nEN.n1003 nEN.n1002 0.0037725
R14634 nEN.n1045 nEN.n1044 0.0037725
R14635 nEN.n1114 nEN.n193 0.00374762
R14636 nEN.n759 nEN.n758 0.0037285
R14637 nEN.n49 nEN.n48 0.0037285
R14638 nEN.n820 nEN.n819 0.00370639
R14639 nEN.n1338 nEN.n1337 0.00370639
R14640 nEN.n1125 nEN.n1124 0.00369524
R14641 nEN.n1180 nEN.n1179 0.00366216
R14642 nEN.n1261 nEN.n1260 0.00366216
R14643 nEN.n1116 nEN.n196 0.00366216
R14644 nEN.n1111 nEN.n1110 0.00364005
R14645 nEN.n329 nEN.n328 0.00363514
R14646 nEN.n389 nEN.n364 0.00363514
R14647 nEN.n1151 nEN.n1150 0.00363514
R14648 nEN.n1291 nEN.n1290 0.00363514
R14649 nEN.n850 nEN.n721 0.00359048
R14650 nEN.n998 nEN.n252 0.00358532
R14651 nEN.n1018 nEN.n1015 0.00358218
R14652 nEN.n316 nEN.n315 0.00357902
R14653 nEN.n379 nEN.n378 0.00357902
R14654 nEN.n941 nEN.n940 0.00357098
R14655 nEN.n1042 nEN.n1041 0.00357098
R14656 nEN.n1188 nEN.n1187 0.00348526
R14657 nEN.n1253 nEN.n1252 0.00348526
R14658 nEN.n965 nEN.n964 0.003457
R14659 nEN.n1068 nEN.n1067 0.003457
R14660 nEN.n263 nEN.n259 0.00344926
R14661 nEN.n212 nEN.n207 0.00344926
R14662 nEN.n833 nEN.n739 0.00344103
R14663 nEN.n816 nEN.n815 0.00344103
R14664 nEN.n1351 nEN.n29 0.00344103
R14665 nEN.n1334 nEN.n1333 0.00344103
R14666 nEN.n990 nEN.n256 0.00343273
R14667 nEN.n1097 nEN.n1096 0.00343273
R14668 nEN.n957 nEN.n956 0.00341839
R14669 nEN.n220 nEN.n219 0.00341839
R14670 nEN.n1062 nEN.n222 0.00341837
R14671 nEN.n954 nEN.n278 0.00341837
R14672 nEN.n849 nEN.n848 0.00335476
R14673 nEN.n1163 nEN.n163 0.00335258
R14674 nEN.n1285 nEN.n1284 0.00335258
R14675 nEN.n956 nEN.n276 0.0033136
R14676 nEN.n1055 nEN.n220 0.0033136
R14677 nEN.n433 nEN.n347 0.00331081
R14678 nEN.n590 nEN.n422 0.00331081
R14679 nEN.n1210 nEN.n1209 0.00331081
R14680 nEN.n1230 nEN.n130 0.00331081
R14681 nEN.n726 nEN.n370 0.00331081
R14682 nEN.n16 nEN.n9 0.00331081
R14683 nEN.n925 nEN.n289 0.00331081
R14684 nEN.n1033 nEN.n1032 0.00331081
R14685 nEN.n266 nEN.n259 0.00330444
R14686 nEN.n1080 nEN.n207 0.00330444
R14687 nEN.n993 nEN.n256 0.0032992
R14688 nEN.n1096 nEN.n1095 0.0032992
R14689 nEN.n964 nEN.n963 0.00329663
R14690 nEN.n1069 nEN.n1068 0.00329663
R14691 nEN.n1122 nEN.n194 0.00324201
R14692 nEN.n1207 nEN.n1206 0.00319779
R14693 nEN.n1236 nEN.n127 0.00319779
R14694 nEN.n804 nEN.n803 0.00319779
R14695 nEN.n1322 nEN.n1321 0.00319779
R14696 nEN.n1123 nEN.n192 0.00319779
R14697 nEN.n846 nEN.n724 0.00317568
R14698 nEN.n1364 nEN.n14 0.00317568
R14699 nEN.n932 nEN.n931 0.00317568
R14700 nEN.n1039 nEN.n233 0.00317568
R14701 nEN.n940 nEN.n939 0.00316007
R14702 nEN.n1043 nEN.n1042 0.00316007
R14703 nEN.n1001 nEN.n252 0.00314581
R14704 nEN.n851 nEN.n371 0.00310934
R14705 nEN.n828 nEN.n740 0.00309459
R14706 nEN.n1346 nEN.n30 0.00309459
R14707 nEN.n960 nEN.n959 0.00309459
R14708 nEN.n1073 nEN.n1072 0.00309459
R14709 nEN.n1144 nEN.n1143 0.003043
R14710 nEN.n1307 nEN.n1306 0.003043
R14711 nEN.n478 nEN.n476 0.0029881
R14712 nEN.n513 nEN.n512 0.0029881
R14713 nEN.n528 nEN.n447 0.0029881
R14714 nEN.n630 nEN.n629 0.0029881
R14715 nEN.n939 nEN.n938 0.00298054
R14716 nEN.n1002 nEN.n1001 0.00298054
R14717 nEN.n1044 nEN.n1043 0.00298054
R14718 nEN.n645 nEN.n404 0.0029619
R14719 nEN.n679 nEN.n678 0.0029619
R14720 nEN.n266 nEN.n260 0.00293083
R14721 nEN.n1080 nEN.n209 0.00293083
R14722 nEN.n963 nEN.n962 0.0029237
R14723 nEN.n1070 nEN.n1069 0.0029237
R14724 nEN.n1213 nEN.n138 0.00291032
R14725 nEN.n1217 nEN.n1216 0.00291032
R14726 nEN.n722 nEN.n372 0.00291032
R14727 nEN.n794 nEN.n786 0.00291032
R14728 nEN.n1367 nEN.n11 0.00291032
R14729 nEN.n91 nEN.n75 0.00291032
R14730 nEN.n1013 nEN.n245 0.00291032
R14731 nEN.n191 nEN.n190 0.00291032
R14732 nEN.n957 nEN.n274 0.00289527
R14733 nEN.n990 nEN.n989 0.00289527
R14734 nEN.n1064 nEN.n219 0.00289527
R14735 nEN.n1097 nEN.n206 0.00289527
R14736 nEN.n316 nEN.n307 0.00287188
R14737 nEN.n715 nEN.n379 0.00284569
R14738 nEN.n249 nEN.n246 0.00283826
R14739 nEN.n1311 nEN.n95 0.00283095
R14740 nEN.n294 nEN.n291 0.00279542
R14741 nEN.n237 nEN.n234 0.00279542
R14742 nEN.n280 nEN.n277 0.00276679
R14743 nEN.n224 nEN.n221 0.00276679
R14744 nEN.n174 nEN.n173 0.00275553
R14745 nEN.n1288 nEN.n104 0.00275553
R14746 nEN.n183 nEN.n181 0.00273342
R14747 nEN.n1313 nEN.n90 0.00273342
R14748 nEN.n318 nEN.n307 0.00272619
R14749 nEN.n319 nEN.n318 0.00272619
R14750 nEN.n913 nEN.n912 0.00272619
R14751 nEN.n911 nEN.n325 0.00272619
R14752 nEN.n902 nEN.n901 0.00272619
R14753 nEN.n470 nEN.n467 0.00272619
R14754 nEN.n475 nEN.n467 0.00272619
R14755 nEN.n477 nEN.n463 0.00272619
R14756 nEN.n485 nEN.n463 0.00272619
R14757 nEN.n493 nEN.n460 0.00272619
R14758 nEN.n494 nEN.n493 0.00272619
R14759 nEN.n503 nEN.n502 0.00272619
R14760 nEN.n504 nEN.n503 0.00272619
R14761 nEN.n514 nEN.n454 0.00272619
R14762 nEN.n518 nEN.n454 0.00272619
R14763 nEN.n526 nEN.n450 0.00272619
R14764 nEN.n527 nEN.n526 0.00272619
R14765 nEN.n535 nEN.n534 0.00272619
R14766 nEN.n536 nEN.n444 0.00272619
R14767 nEN.n548 nEN.n442 0.00272619
R14768 nEN.n560 nEN.n438 0.00272619
R14769 nEN.n561 nEN.n560 0.00272619
R14770 nEN.n567 nEN.n566 0.00272619
R14771 nEN.n569 nEN.n567 0.00272619
R14772 nEN.n569 nEN.n568 0.00272619
R14773 nEN.n578 nEN.n577 0.00272619
R14774 nEN.n587 nEN.n586 0.00272619
R14775 nEN.n586 nEN.n424 0.00272619
R14776 nEN.n596 nEN.n595 0.00272619
R14777 nEN.n595 nEN.n420 0.00272619
R14778 nEN.n602 nEN.n420 0.00272619
R14779 nEN.n610 nEN.n417 0.00272619
R14780 nEN.n611 nEN.n610 0.00272619
R14781 nEN.n620 nEN.n619 0.00272619
R14782 nEN.n621 nEN.n620 0.00272619
R14783 nEN.n635 nEN.n411 0.00272619
R14784 nEN.n644 nEN.n643 0.00272619
R14785 nEN.n652 nEN.n651 0.00272619
R14786 nEN.n653 nEN.n401 0.00272619
R14787 nEN.n665 nEN.n399 0.00272619
R14788 nEN.n677 nEN.n395 0.00272619
R14789 nEN.n678 nEN.n677 0.00272619
R14790 nEN.n685 nEN.n393 0.00272619
R14791 nEN.n686 nEN.n685 0.00272619
R14792 nEN.n687 nEN.n686 0.00272619
R14793 nEN.n695 nEN.n694 0.00272619
R14794 nEN.n695 nEN.n387 0.00272619
R14795 nEN.n704 nEN.n385 0.00272619
R14796 nEN.n705 nEN.n704 0.00272619
R14797 nEN.n714 nEN.n713 0.00272619
R14798 nEN.n716 nEN.n715 0.00272619
R14799 nEN.n319 nEN.n304 0.0027
R14800 nEN.n912 nEN.n911 0.0027
R14801 nEN.n902 nEN.n327 0.0027
R14802 nEN.n470 nEN.n469 0.0027
R14803 nEN.n478 nEN.n477 0.0027
R14804 nEN.n504 nEN.n456 0.0027
R14805 nEN.n536 nEN.n535 0.0027
R14806 nEN.n544 nEN.n442 0.0027
R14807 nEN.n550 nEN.n438 0.0027
R14808 nEN.n578 nEN.n576 0.0027
R14809 nEN.n587 nEN.n585 0.0027
R14810 nEN.n621 nEN.n413 0.0027
R14811 nEN.n631 nEN.n411 0.0027
R14812 nEN.n643 nEN.n407 0.0027
R14813 nEN.n653 nEN.n652 0.0027
R14814 nEN.n661 nEN.n399 0.0027
R14815 nEN.n667 nEN.n395 0.0027
R14816 nEN.n707 nEN.n705 0.0027
R14817 nEN.n716 nEN.n714 0.0027
R14818 nEN.n512 nEN.n456 0.00264762
R14819 nEN.n651 nEN.n404 0.00264762
R14820 nEN.n834 nEN.n737 0.00264496
R14821 nEN.n1352 nEN.n27 0.00264496
R14822 nEN.n781 nEN.n764 0.00262285
R14823 nEN.n70 nEN.n54 0.00262285
R14824 nEN.n994 nEN.n254 0.00262285
R14825 nEN.n1094 nEN.n1091 0.00262285
R14826 nEN.n528 nEN.n527 0.00262143
R14827 nEN.n631 nEN.n630 0.00262143
R14828 nEN.n151 nEN.n148 0.00260074
R14829 nEN.n1240 nEN.n117 0.00260074
R14830 nEN.n480 nEN.n466 0.00257862
R14831 nEN.n680 nEN.n394 0.00257862
R14832 nEN.n629 nEN.n413 0.00256905
R14833 nEN.n524 nEN.n342 0.00255405
R14834 nEN.n625 nEN.n409 0.00255405
R14835 nEN.n1185 nEN.n1184 0.00255405
R14836 nEN.n1250 nEN.n116 0.00255405
R14837 nEN.n1374 nEN.n4 0.00255405
R14838 nEN.n534 nEN.n447 0.00254286
R14839 nEN.n645 nEN.n644 0.00254286
R14840 nEN.n530 nEN.n448 0.0025344
R14841 nEN.n514 nEN.n513 0.00251667
R14842 nEN.n628 nEN.n627 0.00251228
R14843 nEN.n1019 nEN.n1018 0.00249519
R14844 nEN.n313 nEN.n312 0.0024936
R14845 nEN.n476 nEN.n475 0.00246429
R14846 nEN.n679 nEN.n393 0.00246429
R14847 nEN.n1167 nEN.n153 0.00244595
R14848 nEN.n1264 nEN.n113 0.00244595
R14849 nEN.n495 nEN.n494 0.0024381
R14850 nEN.n661 nEN.n660 0.0024381
R14851 nEN.n511 nEN.n510 0.00242383
R14852 nEN.n647 nEN.n405 0.00242383
R14853 nEN.n1115 nEN.n1114 0.00238571
R14854 nEN.n721 nEN.n720 0.00238571
R14855 nEN.n907 nEN.n906 0.00238571
R14856 nEN.n900 nEN.n332 0.00238571
R14857 nEN.n487 nEN.n486 0.00238571
R14858 nEN.n495 nEN.n458 0.00238571
R14859 nEN.n520 nEN.n519 0.00238571
R14860 nEN.n543 nEN.n542 0.00238571
R14861 nEN.n551 nEN.n549 0.00238571
R14862 nEN.n575 nEN.n431 0.00238571
R14863 nEN.n584 nEN.n427 0.00238571
R14864 nEN.n593 nEN.n424 0.00238571
R14865 nEN.n604 nEN.n603 0.00238571
R14866 nEN.n612 nEN.n415 0.00238571
R14867 nEN.n637 nEN.n636 0.00238571
R14868 nEN.n660 nEN.n659 0.00238571
R14869 nEN.n668 nEN.n666 0.00238571
R14870 nEN.n693 nEN.n391 0.00238571
R14871 nEN.n700 nEN.n699 0.00238571
R14872 nEN.n914 nEN.n303 0.00237961
R14873 nEN.n910 nEN.n909 0.00237961
R14874 nEN.n903 nEN.n331 0.00237961
R14875 nEN.n472 nEN.n471 0.00237961
R14876 nEN.n474 nEN.n472 0.00237961
R14877 nEN.n483 nEN.n464 0.00237961
R14878 nEN.n484 nEN.n483 0.00237961
R14879 nEN.n492 nEN.n461 0.00237961
R14880 nEN.n492 nEN.n459 0.00237961
R14881 nEN.n501 nEN.n457 0.00237961
R14882 nEN.n505 nEN.n457 0.00237961
R14883 nEN.n516 nEN.n515 0.00237961
R14884 nEN.n517 nEN.n516 0.00237961
R14885 nEN.n525 nEN.n451 0.00237961
R14886 nEN.n525 nEN.n449 0.00237961
R14887 nEN.n533 nEN.n446 0.00237961
R14888 nEN.n537 nEN.n445 0.00237961
R14889 nEN.n547 nEN.n546 0.00237961
R14890 nEN.n559 nEN.n558 0.00237961
R14891 nEN.n559 nEN.n437 0.00237961
R14892 nEN.n565 nEN.n434 0.00237961
R14893 nEN.n570 nEN.n434 0.00237961
R14894 nEN.n570 nEN.n435 0.00237961
R14895 nEN.n579 nEN.n430 0.00237961
R14896 nEN.n588 nEN.n425 0.00237961
R14897 nEN.n591 nEN.n425 0.00237961
R14898 nEN.n597 nEN.n421 0.00237961
R14899 nEN.n600 nEN.n421 0.00237961
R14900 nEN.n601 nEN.n600 0.00237961
R14901 nEN.n609 nEN.n418 0.00237961
R14902 nEN.n609 nEN.n416 0.00237961
R14903 nEN.n618 nEN.n414 0.00237961
R14904 nEN.n622 nEN.n414 0.00237961
R14905 nEN.n634 nEN.n633 0.00237961
R14906 nEN.n642 nEN.n406 0.00237961
R14907 nEN.n650 nEN.n403 0.00237961
R14908 nEN.n654 nEN.n402 0.00237961
R14909 nEN.n664 nEN.n663 0.00237961
R14910 nEN.n676 nEN.n675 0.00237961
R14911 nEN.n676 nEN.n394 0.00237961
R14912 nEN.n684 nEN.n683 0.00237961
R14913 nEN.n684 nEN.n392 0.00237961
R14914 nEN.n688 nEN.n392 0.00237961
R14915 nEN.n696 nEN.n388 0.00237961
R14916 nEN.n697 nEN.n696 0.00237961
R14917 nEN.n703 nEN.n702 0.00237961
R14918 nEN.n703 nEN.n383 0.00237961
R14919 nEN.n712 nEN.n376 0.00237961
R14920 nEN.n757 nEN.n753 0.00237961
R14921 nEN.n821 nEN.n753 0.00237961
R14922 nEN.n47 nEN.n43 0.00237961
R14923 nEN.n1339 nEN.n43 0.00237961
R14924 nEN.n311 nEN.n306 0.00237961
R14925 nEN.n927 nEN.n926 0.00237961
R14926 nEN.n984 nEN.n262 0.00237961
R14927 nEN.n984 nEN.n983 0.00237961
R14928 nEN.n1009 nEN.n1008 0.00237961
R14929 nEN.n1035 nEN.n1034 0.00237961
R14930 nEN.n1086 nEN.n211 0.00237961
R14931 nEN.n1086 nEN.n1085 0.00237961
R14932 nEN.n544 nEN.n543 0.00235952
R14933 nEN.n566 nEN.n436 0.00235952
R14934 nEN.n321 nEN.n320 0.00235749
R14935 nEN.n910 nEN.n303 0.00235749
R14936 nEN.n904 nEN.n903 0.00235749
R14937 nEN.n471 nEN.n468 0.00235749
R14938 nEN.n479 nEN.n464 0.00235749
R14939 nEN.n506 nEN.n505 0.00235749
R14940 nEN.n537 nEN.n446 0.00235749
R14941 nEN.n546 nEN.n545 0.00235749
R14942 nEN.n558 nEN.n439 0.00235749
R14943 nEN.n579 nEN.n429 0.00235749
R14944 nEN.n588 nEN.n426 0.00235749
R14945 nEN.n623 nEN.n622 0.00235749
R14946 nEN.n633 nEN.n632 0.00235749
R14947 nEN.n642 nEN.n408 0.00235749
R14948 nEN.n654 nEN.n403 0.00235749
R14949 nEN.n663 nEN.n662 0.00235749
R14950 nEN.n675 nEN.n396 0.00235749
R14951 nEN.n708 nEN.n383 0.00235749
R14952 nEN.n952 nEN.n951 0.00235749
R14953 nEN.n1060 nEN.n1059 0.00235749
R14954 nEN.n612 nEN.n611 0.00233333
R14955 nEN.n511 nEN.n506 0.00231327
R14956 nEN.n650 nEN.n405 0.00231327
R14957 nEN.n323 nEN.n304 0.00230714
R14958 nEN.n707 nEN.n706 0.00230714
R14959 nEN.n713 nEN.n380 0.00230714
R14960 nEN.n529 nEN.n449 0.00229115
R14961 nEN.n632 nEN.n412 0.00229115
R14962 nEN.n1168 nEN.n1167 0.00229115
R14963 nEN.n1271 nEN.n1264 0.00229115
R14964 nEN.n913 nEN.n324 0.00228095
R14965 nEN.n901 nEN.n900 0.00228095
R14966 nEN.n694 nEN.n693 0.00225476
R14967 nEN.n628 nEN.n623 0.00224693
R14968 nEN.n2 nEN 0.0022301
R14969 nEN.n844 nEN.n843 0.00222973
R14970 nEN.n1362 nEN.n1361 0.00222973
R14971 nEN.n935 nEN.n934 0.00222973
R14972 nEN.n1047 nEN.n230 0.00222973
R14973 nEN.n533 nEN.n448 0.00222482
R14974 nEN.n646 nEN.n406 0.00222482
R14975 nEN.n515 nEN.n455 0.0022027
R14976 nEN.n562 nEN.n561 0.00220238
R14977 nEN.n596 nEN.n594 0.00220238
R14978 nEN.n576 nEN.n575 0.00217619
R14979 nEN.n577 nEN.n427 0.00217619
R14980 nEN.n1015 nEN.n1014 0.00217613
R14981 nEN.n474 nEN.n466 0.00215848
R14982 nEN.n683 nEN.n680 0.00215848
R14983 nEN.n496 nEN.n459 0.00213636
R14984 nEN.n662 nEN.n400 0.00213636
R14985 nEN.n1194 nEN.n148 0.00213636
R14986 nEN.n1241 nEN.n1240 0.00213636
R14987 nEN.n782 nEN.n781 0.00211425
R14988 nEN.n71 nEN.n70 0.00211425
R14989 nEN.n997 nEN.n254 0.00211425
R14990 nEN.n1091 nEN.n198 0.00211425
R14991 nEN.n850 nEN.n849 0.00209762
R14992 nEN.n906 nEN.n327 0.00209762
R14993 nEN.n592 nEN.n591 0.00209214
R14994 nEN.n837 nEN.n737 0.00209214
R14995 nEN.n1355 nEN.n27 0.00209214
R14996 nEN.n953 nEN.n280 0.00209214
R14997 nEN.n1061 nEN.n224 0.00209214
R14998 nEN.n699 nEN.n387 0.00207143
R14999 nEN.n545 nEN.n443 0.00207002
R15000 nEN.n565 nEN.n564 0.00207002
R15001 nEN.n613 nEN.n416 0.00204791
R15002 nEN.n322 nEN.n321 0.0020258
R15003 nEN.n708 nEN.n384 0.0020258
R15004 nEN.n712 nEN.n381 0.0020258
R15005 nEN.n549 nEN.n548 0.00201905
R15006 nEN.n832 nEN.n738 0.00201351
R15007 nEN.n1350 nEN.n28 0.00201351
R15008 nEN.n949 nEN.n275 0.00201351
R15009 nEN.n1057 nEN.n1056 0.00201351
R15010 nEN.n914 nEN.n302 0.00200369
R15011 nEN.n899 nEN.n331 0.00200369
R15012 nEN.n175 nEN.n174 0.00200369
R15013 nEN.n1289 nEN.n1288 0.00200369
R15014 nEN.n719 nEN.n375 0.00200107
R15015 nEN.n314 nEN.n313 0.00200107
R15016 nEN.n312 nEN.n293 0.00200107
R15017 nEN.n604 nEN.n417 0.00199286
R15018 nEN.n692 nEN.n388 0.00198157
R15019 nEN.n563 nEN.n437 0.00193735
R15020 nEN.n597 nEN.n423 0.00193735
R15021 nEN.n574 nEN.n429 0.00191523
R15022 nEN.n430 nEN.n428 0.00191523
R15023 nEN.n718 nEN.n717 0.00191523
R15024 nEN.n1313 nEN.n94 0.00191523
R15025 nEN.n317 nEN.n306 0.00191523
R15026 nEN.n311 nEN.n310 0.00191523
R15027 nEN.n487 nEN.n460 0.00191429
R15028 nEN.n666 nEN.n665 0.00191429
R15029 nEN.n500 nEN.n499 0.00187101
R15030 nEN.n951 nEN.n281 0.00185493
R15031 nEN.n1059 nEN.n225 0.00185493
R15032 nEN.n905 nEN.n904 0.00184889
R15033 nEN.n658 nEN.n657 0.00184889
R15034 nEN.n1213 nEN.n1212 0.00184889
R15035 nEN.n1220 nEN.n1217 0.00184889
R15036 nEN.n851 nEN.n372 0.00184889
R15037 nEN.n798 nEN.n794 0.00184889
R15038 nEN.n1368 nEN.n1367 0.00184889
R15039 nEN.n92 nEN.n91 0.00184889
R15040 nEN.n928 nEN.n294 0.00184889
R15041 nEN.n1021 nEN.n1013 0.00184889
R15042 nEN.n1036 nEN.n237 0.00184889
R15043 nEN.n1131 nEN.n190 0.00184889
R15044 nEN.n637 nEN.n407 0.00183571
R15045 nEN.n698 nEN.n697 0.00182678
R15046 nEN.n519 nEN.n518 0.00180952
R15047 nEN.n508 nEN.n452 0.0017973
R15048 nEN.n641 nEN.n357 0.0017973
R15049 nEN.n1177 nEN.n152 0.0017973
R15050 nEN.n1258 nEN.n1257 0.0017973
R15051 nEN.n926 nEN.n290 0.0017897
R15052 nEN.n1034 nEN.n238 0.0017897
R15053 nEN.n541 nEN.n540 0.00178256
R15054 nEN.n547 nEN.n441 0.00178256
R15055 nEN.n617 nEN.n616 0.00178256
R15056 nEN.n605 nEN.n418 0.00176044
R15057 nEN.n1124 nEN.n193 0.00175714
R15058 nEN.n520 nEN.n450 0.00173095
R15059 nEN.n636 nEN.n635 0.00173095
R15060 nEN.n898 nEN.n333 0.00171622
R15061 nEN.n1008 nEN.n250 0.00171347
R15062 nEN.n488 nEN.n461 0.0016941
R15063 nEN.n664 nEN.n398 0.0016941
R15064 nEN.n691 nEN.n689 0.0016941
R15065 nEN.n1144 nEN.n172 0.0016941
R15066 nEN.n1307 nEN.n97 0.0016941
R15067 nEN.n668 nEN.n667 0.00165238
R15068 nEN.n573 nEN.n432 0.00162776
R15069 nEN.n583 nEN.n582 0.00162776
R15070 nEN.n638 nEN.n408 0.00162776
R15071 nEN.n373 nEN.n371 0.00162776
R15072 nEN.n486 nEN.n485 0.00162619
R15073 nEN.n517 nEN.n453 0.00160565
R15074 nEN.n846 nEN.n845 0.00158354
R15075 nEN.n1364 nEN.n1363 0.00158354
R15076 nEN.n931 nEN.n288 0.00158354
R15077 nEN.n1040 nEN.n1039 0.00158354
R15078 nEN.n908 nEN.n326 0.00156143
R15079 nEN.n701 nEN.n386 0.00156143
R15080 nEN.n1206 nEN.n1205 0.00156143
R15081 nEN.n1236 nEN.n1235 0.00156143
R15082 nEN.n804 nEN.n785 0.00156143
R15083 nEN.n1322 nEN.n74 0.00156143
R15084 nEN.n1010 nEN.n249 0.00156143
R15085 nEN.n1123 nEN.n1122 0.00156143
R15086 nEN.n551 nEN.n550 0.00154762
R15087 nEN.n603 nEN.n602 0.00154762
R15088 nEN.n521 nEN.n451 0.00153931
R15089 nEN.n634 nEN.n410 0.00153931
R15090 nEN.n553 nEN.n552 0.00149509
R15091 nEN.n1117 nEN.n194 0.00149509
R15092 nEN.n606 nEN.n419 0.00147297
R15093 nEN.n669 nEN.n396 0.00147297
R15094 nEN.n907 nEN.n325 0.00146905
R15095 nEN.n700 nEN.n385 0.00146905
R15096 nEN.n484 nEN.n462 0.00145086
R15097 nEN.n489 nEN.n462 0.00140663
R15098 nEN.n670 nEN.n669 0.00140663
R15099 nEN.n1163 nEN.n1162 0.00140663
R15100 nEN.n1285 nEN.n106 0.00140663
R15101 nEN.n585 nEN.n584 0.00139048
R15102 nEN.n552 nEN.n439 0.00138452
R15103 nEN.n601 nEN.n419 0.00138452
R15104 nEN.n324 nEN.n323 0.00136429
R15105 nEN.n562 nEN.n436 0.00136429
R15106 nEN.n568 nEN.n431 0.00136429
R15107 nEN.n522 nEN.n521 0.00134029
R15108 nEN.n639 nEN.n410 0.00134029
R15109 nEN.n594 nEN.n593 0.00133809
R15110 nEN.n706 nEN.n380 0.00133809
R15111 nEN.n909 nEN.n908 0.00131818
R15112 nEN.n702 nEN.n701 0.00131818
R15113 nEN.n1010 nEN.n1009 0.00131818
R15114 nEN.n830 nEN.n739 0.00129607
R15115 nEN.n816 nEN.n763 0.00129607
R15116 nEN.n1348 nEN.n29 0.00129607
R15117 nEN.n1334 nEN.n53 0.00129607
R15118 nEN.n469 nEN.n332 0.00128571
R15119 nEN.n687 nEN.n391 0.00128571
R15120 nEN.n522 nEN.n453 0.00125184
R15121 nEN.n583 nEN.n426 0.00125184
R15122 nEN.n639 nEN.n638 0.00125184
R15123 nEN.n1188 nEN.n150 0.00125184
R15124 nEN.n1254 nEN.n1253 0.00125184
R15125 nEN.n322 nEN.n302 0.00122973
R15126 nEN.n564 nEN.n563 0.00122973
R15127 nEN.n435 nEN.n432 0.00122973
R15128 nEN.n592 nEN.n423 0.00120762
R15129 nEN.n384 nEN.n381 0.00120762
R15130 nEN.n542 nEN.n444 0.00120714
R15131 nEN.n619 nEN.n415 0.00120714
R15132 nEN.n489 nEN.n488 0.0011855
R15133 nEN.n670 nEN.n398 0.0011855
R15134 nEN.n468 nEN.n333 0.00116339
R15135 nEN.n689 nEN.n688 0.00116339
R15136 nEN.n840 nEN.n733 0.00114865
R15137 nEN.n1358 nEN.n23 0.00114865
R15138 nEN.n943 nEN.n286 0.00114865
R15139 nEN.n232 nEN.n231 0.00114865
R15140 nEN.n659 nEN.n401 0.00112857
R15141 nEN.n606 nEN.n605 0.00111916
R15142 nEN.n502 nEN.n458 0.00110238
R15143 nEN.n541 nEN.n445 0.00109705
R15144 nEN.n553 nEN.n441 0.00109705
R15145 nEN.n618 nEN.n617 0.00109705
R15146 nEN.n1181 nEN.n1180 0.00109705
R15147 nEN.n1261 nEN.n115 0.00109705
R15148 nEN.n1117 nEN.n1116 0.00109705
R15149 nEN.n819 nEN.n754 0.00105283
R15150 nEN.n1337 nEN.n44 0.00105283
R15151 nEN.n1310 nEN.n94 0.00105283
R15152 nEN.n572 nEN.n348 0.00104054
R15153 nEN.n1224 nEN.n134 0.00104054
R15154 nEN.n905 nEN.n326 0.00103071
R15155 nEN.n658 nEN.n402 0.00103071
R15156 nEN.n698 nEN.n386 0.00103071
R15157 nEN.n717 nEN.n377 0.00103071
R15158 nEN.n759 nEN.n741 0.00103071
R15159 nEN.n49 nEN.n31 0.00103071
R15160 nEN.n317 nEN.n308 0.00103071
R15161 nEN.n928 nEN.n927 0.00103071
R15162 nEN.n1036 nEN.n1035 0.00103071
R15163 nEN.n501 nEN.n500 0.0010086
R15164 nEN.n574 nEN.n573 0.000964373
R15165 nEN.n582 nEN.n428 0.000964373
R15166 nEN.n374 nEN.n373 0.000964373
R15167 nEN.n310 nEN.n309 0.000964373
R15168 nEN.n1130 nEN.n1129 0.000964373
R15169 nEN.n164 nEN.n161 0.00094226
R15170 nEN.n1269 nEN.n1268 0.00094226
R15171 nEN.n836 nEN.n734 0.000932432
R15172 nEN.n1354 nEN.n24 0.000932432
R15173 nEN.n287 nEN.n282 0.000932432
R15174 nEN.n1054 nEN.n1053 0.000932432
R15175 nEN.n320 nEN.n306 0.000898034
R15176 nEN.n692 nEN.n691 0.000898034
R15177 nEN.n899 nEN.n898 0.000875921
R15178 nEN.n718 nEN.n376 0.000853808
R15179 nEN.n1110 nEN.n1109 0.000831695
R15180 nEN.n1113 nEN.n1112 0.000814286
R15181 nEN.n540 nEN.n443 0.000809582
R15182 nEN.n616 nEN.n613 0.000809582
R15183 nEN.n1192 nEN.n140 0.000787469
R15184 nEN.n128 nEN.n125 0.000787469
R15185 nEN.n953 nEN.n952 0.000787469
R15186 nEN.n1061 nEN.n1060 0.000787469
R15187 nEN.n736 nEN.n735 0.000765356
R15188 nEN.n807 nEN.n783 0.000765356
R15189 nEN.n26 nEN.n25 0.000765356
R15190 nEN.n1325 nEN.n72 0.000765356
R15191 nEN.n1111 nEN.n196 0.000765356
R15192 nEN.n657 nEN.n400 0.000743243
R15193 nEN.n499 nEN.n496 0.00072113
R15194 nEN.n897 nEN.n896 0.000716216
R15195 nEN.n690 nEN.n363 0.000716216
R15196 nEN.n178 nEN.n177 0.000716216
R15197 nEN.n1297 nEN.n1296 0.000716216
R15198 nEN.n510 nEN.n455 0.000676904
R15199 nEN.n647 nEN.n646 0.000654791
R15200 nEN.n1148 nEN.n1147 0.000654791
R15201 nEN.n1294 nEN.n1293 0.000654791
R15202 nEN.n627 nEN.n412 0.000588452
R15203 nEN.n530 nEN.n529 0.000566339
R15204 nEN.n480 nEN.n479 0.000522113
R15205 nEN.n184 nEN.n183 0.000522113
R15206 CLK_IN.n6 CLK_IN.n0 28.593
R15207 CLK_IN.n1384 CLK_IN 23.8353
R15208 CLK_IN.n3 CLK_IN.n2 17.8375
R15209 CLK_IN.n5 CLK_IN.n4 16.216
R15210 CLK_IN.n9 CLK_IN.n8 15.8163
R15211 CLK_IN.n9 CLK_IN.n7 15.6165
R15212 CLK_IN.n3 CLK_IN.n1 15.2022
R15213 CLK_IN.n6 CLK_IN.n5 9.0115
R15214 CLK_IN.n10 CLK_IN.n9 9.0005
R15215 CLK_IN.n867 CLK_IN.n866 2.2505
R15216 CLK_IN.n873 CLK_IN.n872 2.2505
R15217 CLK_IN.n888 CLK_IN.n219 2.2505
R15218 CLK_IN.n221 CLK_IN.n217 2.2505
R15219 CLK_IN.n937 CLK_IN.n201 2.2505
R15220 CLK_IN.n945 CLK_IN.n199 2.2505
R15221 CLK_IN.n974 CLK_IN.n13 2.2505
R15222 CLK_IN.n1380 CLK_IN.n15 2.2505
R15223 CLK_IN.n1379 CLK_IN.n16 2.2505
R15224 CLK_IN.n1375 CLK_IN.n19 2.2505
R15225 CLK_IN.n1373 CLK_IN.n21 2.2505
R15226 CLK_IN.n1369 CLK_IN.n24 2.2505
R15227 CLK_IN.n1367 CLK_IN.n26 2.2505
R15228 CLK_IN.n1363 CLK_IN.n29 2.2505
R15229 CLK_IN.n1361 CLK_IN.n31 2.2505
R15230 CLK_IN.n88 CLK_IN.n76 2.2505
R15231 CLK_IN.n500 CLK_IN.n79 2.2505
R15232 CLK_IN.n654 CLK_IN.n495 2.2505
R15233 CLK_IN.n658 CLK_IN.n492 2.2505
R15234 CLK_IN.n660 CLK_IN.n490 2.2505
R15235 CLK_IN.n664 CLK_IN.n487 2.2505
R15236 CLK_IN.n666 CLK_IN.n485 2.2505
R15237 CLK_IN.n518 CLK_IN.n483 2.2505
R15238 CLK_IN.n671 CLK_IN.n481 2.2505
R15239 CLK_IN.n580 CLK_IN.n478 2.2505
R15240 CLK_IN.n677 CLK_IN.n476 2.2505
R15241 CLK_IN.n556 CLK_IN.n473 2.2505
R15242 CLK_IN.n683 CLK_IN.n471 2.2505
R15243 CLK_IN.n534 CLK_IN.n466 2.2505
R15244 CLK_IN.n465 CLK_IN.n464 2.2505
R15245 CLK_IN.n1305 CLK_IN.n76 2.2505
R15246 CLK_IN.n79 CLK_IN.n78 2.2505
R15247 CLK_IN.n655 CLK_IN.n654 2.2505
R15248 CLK_IN.n658 CLK_IN.n657 2.2505
R15249 CLK_IN.n661 CLK_IN.n660 2.2505
R15250 CLK_IN.n664 CLK_IN.n663 2.2505
R15251 CLK_IN.n667 CLK_IN.n666 2.2505
R15252 CLK_IN.n668 CLK_IN.n483 2.2505
R15253 CLK_IN.n671 CLK_IN.n479 2.2505
R15254 CLK_IN.n674 CLK_IN.n478 2.2505
R15255 CLK_IN.n677 CLK_IN.n474 2.2505
R15256 CLK_IN.n680 CLK_IN.n473 2.2505
R15257 CLK_IN.n683 CLK_IN.n469 2.2505
R15258 CLK_IN.n686 CLK_IN.n466 2.2505
R15259 CLK_IN.n468 CLK_IN.n465 2.2505
R15260 CLK_IN.n701 CLK_IN.n450 2.2505
R15261 CLK_IN.n702 CLK_IN.n449 2.2505
R15262 CLK_IN.n448 CLK_IN.n432 2.2505
R15263 CLK_IN.n715 CLK_IN.n431 2.2505
R15264 CLK_IN.n716 CLK_IN.n430 2.2505
R15265 CLK_IN.n429 CLK_IN.n414 2.2505
R15266 CLK_IN.n727 CLK_IN.n413 2.2505
R15267 CLK_IN.n728 CLK_IN.n412 2.2505
R15268 CLK_IN.n411 CLK_IN.n398 2.2505
R15269 CLK_IN.n410 CLK_IN.n409 2.2505
R15270 CLK_IN.n399 CLK_IN.n379 2.2505
R15271 CLK_IN.n741 CLK_IN.n378 2.2505
R15272 CLK_IN.n742 CLK_IN.n377 2.2505
R15273 CLK_IN.n376 CLK_IN.n370 2.2505
R15274 CLK_IN.n375 CLK_IN.n374 2.2505
R15275 CLK_IN.n373 CLK_IN.n372 2.2505
R15276 CLK_IN.n371 CLK_IN.n348 2.2505
R15277 CLK_IN.n765 CLK_IN.n347 2.2505
R15278 CLK_IN.n766 CLK_IN.n346 2.2505
R15279 CLK_IN.n345 CLK_IN.n332 2.2505
R15280 CLK_IN.n779 CLK_IN.n331 2.2505
R15281 CLK_IN.n780 CLK_IN.n330 2.2505
R15282 CLK_IN.n329 CLK_IN.n327 2.2505
R15283 CLK_IN.n328 CLK_IN.n305 2.2505
R15284 CLK_IN.n792 CLK_IN.n304 2.2505
R15285 CLK_IN.n793 CLK_IN.n303 2.2505
R15286 CLK_IN.n302 CLK_IN.n282 2.2505
R15287 CLK_IN.n301 CLK_IN.n300 2.2505
R15288 CLK_IN.n299 CLK_IN.n283 2.2505
R15289 CLK_IN.n298 CLK_IN.n287 2.2505
R15290 CLK_IN.n286 CLK_IN.n284 2.2505
R15291 CLK_IN.n285 CLK_IN.n256 2.2505
R15292 CLK_IN.n819 CLK_IN.n255 2.2505
R15293 CLK_IN.n820 CLK_IN.n254 2.2505
R15294 CLK_IN.n821 CLK_IN.n820 2.2505
R15295 CLK_IN.n819 CLK_IN.n818 2.2505
R15296 CLK_IN.n288 CLK_IN.n256 2.2505
R15297 CLK_IN.n293 CLK_IN.n284 2.2505
R15298 CLK_IN.n298 CLK_IN.n297 2.2505
R15299 CLK_IN.n299 CLK_IN.n275 2.2505
R15300 CLK_IN.n300 CLK_IN.n276 2.2505
R15301 CLK_IN.n282 CLK_IN.n278 2.2505
R15302 CLK_IN.n794 CLK_IN.n793 2.2505
R15303 CLK_IN.n792 CLK_IN.n791 2.2505
R15304 CLK_IN.n321 CLK_IN.n305 2.2505
R15305 CLK_IN.n327 CLK_IN.n326 2.2505
R15306 CLK_IN.n781 CLK_IN.n780 2.2505
R15307 CLK_IN.n779 CLK_IN.n778 2.2505
R15308 CLK_IN.n341 CLK_IN.n332 2.2505
R15309 CLK_IN.n767 CLK_IN.n766 2.2505
R15310 CLK_IN.n765 CLK_IN.n764 2.2505
R15311 CLK_IN.n359 CLK_IN.n348 2.2505
R15312 CLK_IN.n373 CLK_IN.n363 2.2505
R15313 CLK_IN.n374 CLK_IN.n364 2.2505
R15314 CLK_IN.n370 CLK_IN.n366 2.2505
R15315 CLK_IN.n743 CLK_IN.n742 2.2505
R15316 CLK_IN.n741 CLK_IN.n740 2.2505
R15317 CLK_IN.n400 CLK_IN.n379 2.2505
R15318 CLK_IN.n409 CLK_IN.n408 2.2505
R15319 CLK_IN.n398 CLK_IN.n396 2.2505
R15320 CLK_IN.n729 CLK_IN.n728 2.2505
R15321 CLK_IN.n727 CLK_IN.n726 2.2505
R15322 CLK_IN.n426 CLK_IN.n414 2.2505
R15323 CLK_IN.n717 CLK_IN.n716 2.2505
R15324 CLK_IN.n715 CLK_IN.n714 2.2505
R15325 CLK_IN.n444 CLK_IN.n432 2.2505
R15326 CLK_IN.n703 CLK_IN.n702 2.2505
R15327 CLK_IN.n701 CLK_IN.n700 2.2505
R15328 CLK_IN.n1357 CLK_IN.n34 2.2505
R15329 CLK_IN.n1356 CLK_IN.n35 2.2505
R15330 CLK_IN.n1355 CLK_IN.n36 2.2505
R15331 CLK_IN.n1156 CLK_IN.n37 2.2505
R15332 CLK_IN.n1351 CLK_IN.n39 2.2505
R15333 CLK_IN.n1350 CLK_IN.n40 2.2505
R15334 CLK_IN.n1349 CLK_IN.n41 2.2505
R15335 CLK_IN.n1171 CLK_IN.n42 2.2505
R15336 CLK_IN.n1345 CLK_IN.n44 2.2505
R15337 CLK_IN.n1344 CLK_IN.n45 2.2505
R15338 CLK_IN.n1343 CLK_IN.n46 2.2505
R15339 CLK_IN.n114 CLK_IN.n47 2.2505
R15340 CLK_IN.n1339 CLK_IN.n49 2.2505
R15341 CLK_IN.n1338 CLK_IN.n50 2.2505
R15342 CLK_IN.n1337 CLK_IN.n51 2.2505
R15343 CLK_IN.n1210 CLK_IN.n52 2.2505
R15344 CLK_IN.n1333 CLK_IN.n54 2.2505
R15345 CLK_IN.n1332 CLK_IN.n55 2.2505
R15346 CLK_IN.n1331 CLK_IN.n56 2.2505
R15347 CLK_IN.n1228 CLK_IN.n57 2.2505
R15348 CLK_IN.n1327 CLK_IN.n59 2.2505
R15349 CLK_IN.n1326 CLK_IN.n60 2.2505
R15350 CLK_IN.n1325 CLK_IN.n61 2.2505
R15351 CLK_IN.n1245 CLK_IN.n62 2.2505
R15352 CLK_IN.n1321 CLK_IN.n64 2.2505
R15353 CLK_IN.n1320 CLK_IN.n65 2.2505
R15354 CLK_IN.n1319 CLK_IN.n66 2.2505
R15355 CLK_IN.n97 CLK_IN.n67 2.2505
R15356 CLK_IN.n1315 CLK_IN.n69 2.2505
R15357 CLK_IN.n1314 CLK_IN.n70 2.2505
R15358 CLK_IN.n1313 CLK_IN.n71 2.2505
R15359 CLK_IN.n1284 CLK_IN.n72 2.2505
R15360 CLK_IN.n1309 CLK_IN.n74 2.2505
R15361 CLK_IN.n1308 CLK_IN.n75 2.2505
R15362 CLK_IN.n1308 CLK_IN.n73 2.2505
R15363 CLK_IN.n1310 CLK_IN.n1309 2.2505
R15364 CLK_IN.n1311 CLK_IN.n72 2.2505
R15365 CLK_IN.n1313 CLK_IN.n1312 2.2505
R15366 CLK_IN.n1314 CLK_IN.n68 2.2505
R15367 CLK_IN.n1316 CLK_IN.n1315 2.2505
R15368 CLK_IN.n1317 CLK_IN.n67 2.2505
R15369 CLK_IN.n1319 CLK_IN.n1318 2.2505
R15370 CLK_IN.n1320 CLK_IN.n63 2.2505
R15371 CLK_IN.n1322 CLK_IN.n1321 2.2505
R15372 CLK_IN.n1323 CLK_IN.n62 2.2505
R15373 CLK_IN.n1325 CLK_IN.n1324 2.2505
R15374 CLK_IN.n1326 CLK_IN.n58 2.2505
R15375 CLK_IN.n1328 CLK_IN.n1327 2.2505
R15376 CLK_IN.n1329 CLK_IN.n57 2.2505
R15377 CLK_IN.n1331 CLK_IN.n1330 2.2505
R15378 CLK_IN.n1332 CLK_IN.n53 2.2505
R15379 CLK_IN.n1334 CLK_IN.n1333 2.2505
R15380 CLK_IN.n1335 CLK_IN.n52 2.2505
R15381 CLK_IN.n1337 CLK_IN.n1336 2.2505
R15382 CLK_IN.n1338 CLK_IN.n48 2.2505
R15383 CLK_IN.n1340 CLK_IN.n1339 2.2505
R15384 CLK_IN.n1341 CLK_IN.n47 2.2505
R15385 CLK_IN.n1343 CLK_IN.n1342 2.2505
R15386 CLK_IN.n1344 CLK_IN.n43 2.2505
R15387 CLK_IN.n1346 CLK_IN.n1345 2.2505
R15388 CLK_IN.n1347 CLK_IN.n42 2.2505
R15389 CLK_IN.n1349 CLK_IN.n1348 2.2505
R15390 CLK_IN.n1350 CLK_IN.n38 2.2505
R15391 CLK_IN.n1352 CLK_IN.n1351 2.2505
R15392 CLK_IN.n1353 CLK_IN.n37 2.2505
R15393 CLK_IN.n1355 CLK_IN.n1354 2.2505
R15394 CLK_IN.n1356 CLK_IN.n33 2.2505
R15395 CLK_IN.n1358 CLK_IN.n1357 2.2505
R15396 CLK_IN.n868 CLK_IN.n867 2.2505
R15397 CLK_IN.n872 CLK_IN.n871 2.2505
R15398 CLK_IN.n219 CLK_IN.n218 2.2505
R15399 CLK_IN.n915 CLK_IN.n217 2.2505
R15400 CLK_IN.n201 CLK_IN.n200 2.2505
R15401 CLK_IN.n970 CLK_IN.n199 2.2505
R15402 CLK_IN.n13 CLK_IN.n11 2.2505
R15403 CLK_IN.n1380 CLK_IN.n12 2.2505
R15404 CLK_IN.n1379 CLK_IN.n1378 2.2505
R15405 CLK_IN.n1376 CLK_IN.n1375 2.2505
R15406 CLK_IN.n1373 CLK_IN.n1372 2.2505
R15407 CLK_IN.n1370 CLK_IN.n1369 2.2505
R15408 CLK_IN.n1367 CLK_IN.n1366 2.2505
R15409 CLK_IN.n1364 CLK_IN.n1363 2.2505
R15410 CLK_IN.n1361 CLK_IN.n1360 2.2505
R15411 CLK_IN.n1135 CLK_IN.n1134 2.2005
R15412 CLK_IN.n1123 CLK_IN.n1122 2.2005
R15413 CLK_IN.n1121 CLK_IN.n1120 2.2005
R15414 CLK_IN.n1114 CLK_IN.n1113 2.2005
R15415 CLK_IN.n1112 CLK_IN.n1111 2.2005
R15416 CLK_IN.n1105 CLK_IN.n142 2.2005
R15417 CLK_IN.n1096 CLK_IN.n146 2.2005
R15418 CLK_IN.n1098 CLK_IN.n1097 2.2005
R15419 CLK_IN.n1094 CLK_IN.n1093 2.2005
R15420 CLK_IN.n1088 CLK_IN.n149 2.2005
R15421 CLK_IN.n155 CLK_IN.n152 2.2005
R15422 CLK_IN.n1081 CLK_IN.n156 2.2005
R15423 CLK_IN.n1076 CLK_IN.n1075 2.2005
R15424 CLK_IN.n1074 CLK_IN.n1073 2.2005
R15425 CLK_IN.n1068 CLK_IN.n1067 2.2005
R15426 CLK_IN.n1066 CLK_IN.n1065 2.2005
R15427 CLK_IN.n1060 CLK_IN.n1059 2.2005
R15428 CLK_IN.n1058 CLK_IN.n1057 2.2005
R15429 CLK_IN.n1051 CLK_IN.n167 2.2005
R15430 CLK_IN.n1045 CLK_IN.n1044 2.2005
R15431 CLK_IN.n1043 CLK_IN.n1042 2.2005
R15432 CLK_IN.n1033 CLK_IN.n172 2.2005
R15433 CLK_IN.n1035 CLK_IN.n1034 2.2005
R15434 CLK_IN.n1028 CLK_IN.n1027 2.2005
R15435 CLK_IN.n1026 CLK_IN.n1025 2.2005
R15436 CLK_IN.n1019 CLK_IN.n1018 2.2005
R15437 CLK_IN.n1017 CLK_IN.n1016 2.2005
R15438 CLK_IN.n1010 CLK_IN.n1009 2.2005
R15439 CLK_IN.n1008 CLK_IN.n1007 2.2005
R15440 CLK_IN.n1001 CLK_IN.n1000 2.2005
R15441 CLK_IN.n999 CLK_IN.n998 2.2005
R15442 CLK_IN.n992 CLK_IN.n991 2.2005
R15443 CLK_IN.n990 CLK_IN.n989 2.2005
R15444 CLK_IN.n984 CLK_IN.n191 2.2005
R15445 CLK_IN.n975 CLK_IN.n195 2.2005
R15446 CLK_IN.n977 CLK_IN.n976 2.2005
R15447 CLK_IN.n952 CLK_IN.n198 2.2005
R15448 CLK_IN.n947 CLK_IN.n946 2.2005
R15449 CLK_IN.n960 CLK_IN.n203 2.2005
R15450 CLK_IN.n966 CLK_IN.n965 2.2005
R15451 CLK_IN.n941 CLK_IN.n202 2.2005
R15452 CLK_IN.n939 CLK_IN.n938 2.2005
R15453 CLK_IN.n936 CLK_IN.n935 2.2005
R15454 CLK_IN.n928 CLK_IN.n208 2.2005
R15455 CLK_IN.n216 CLK_IN.n212 2.2005
R15456 CLK_IN.n920 CLK_IN.n919 2.2005
R15457 CLK_IN.n903 CLK_IN.n215 2.2005
R15458 CLK_IN.n905 CLK_IN.n222 2.2005
R15459 CLK_IN.n911 CLK_IN.n910 2.2005
R15460 CLK_IN.n896 CLK_IN.n220 2.2005
R15461 CLK_IN.n890 CLK_IN.n889 2.2005
R15462 CLK_IN.n887 CLK_IN.n886 2.2005
R15463 CLK_IN.n881 CLK_IN.n229 2.2005
R15464 CLK_IN.n879 CLK_IN.n233 2.2005
R15465 CLK_IN.n875 CLK_IN.n874 2.2005
R15466 CLK_IN.n848 CLK_IN.n236 2.2005
R15467 CLK_IN.n853 CLK_IN.n844 2.2005
R15468 CLK_IN.n843 CLK_IN.n840 2.2005
R15469 CLK_IN.n860 CLK_IN.n243 2.2005
R15470 CLK_IN.n865 CLK_IN.n864 2.2005
R15471 CLK_IN.n835 CLK_IN.n242 2.2005
R15472 CLK_IN.n90 CLK_IN.n89 2.2005
R15473 CLK_IN.n459 CLK_IN.n453 2.2005
R15474 CLK_IN.n462 CLK_IN.n460 2.2005
R15475 CLK_IN.n691 CLK_IN.n690 2.2005
R15476 CLK_IN.n463 CLK_IN.n461 2.2005
R15477 CLK_IN.n537 CLK_IN.n536 2.2005
R15478 CLK_IN.n539 CLK_IN.n538 2.2005
R15479 CLK_IN.n541 CLK_IN.n540 2.2005
R15480 CLK_IN.n543 CLK_IN.n542 2.2005
R15481 CLK_IN.n545 CLK_IN.n544 2.2005
R15482 CLK_IN.n547 CLK_IN.n546 2.2005
R15483 CLK_IN.n549 CLK_IN.n548 2.2005
R15484 CLK_IN.n551 CLK_IN.n550 2.2005
R15485 CLK_IN.n554 CLK_IN.n553 2.2005
R15486 CLK_IN.n555 CLK_IN.n529 2.2005
R15487 CLK_IN.n559 CLK_IN.n558 2.2005
R15488 CLK_IN.n557 CLK_IN.n527 2.2005
R15489 CLK_IN.n565 CLK_IN.n564 2.2005
R15490 CLK_IN.n566 CLK_IN.n526 2.2005
R15491 CLK_IN.n568 CLK_IN.n567 2.2005
R15492 CLK_IN.n571 CLK_IN.n570 2.2005
R15493 CLK_IN.n573 CLK_IN.n572 2.2005
R15494 CLK_IN.n524 CLK_IN.n523 2.2005
R15495 CLK_IN.n579 CLK_IN.n578 2.2005
R15496 CLK_IN.n581 CLK_IN.n522 2.2005
R15497 CLK_IN.n583 CLK_IN.n582 2.2005
R15498 CLK_IN.n585 CLK_IN.n584 2.2005
R15499 CLK_IN.n587 CLK_IN.n586 2.2005
R15500 CLK_IN.n589 CLK_IN.n588 2.2005
R15501 CLK_IN.n592 CLK_IN.n591 2.2005
R15502 CLK_IN.n590 CLK_IN.n519 2.2005
R15503 CLK_IN.n598 CLK_IN.n597 2.2005
R15504 CLK_IN.n600 CLK_IN.n599 2.2005
R15505 CLK_IN.n602 CLK_IN.n601 2.2005
R15506 CLK_IN.n604 CLK_IN.n603 2.2005
R15507 CLK_IN.n606 CLK_IN.n605 2.2005
R15508 CLK_IN.n608 CLK_IN.n607 2.2005
R15509 CLK_IN.n610 CLK_IN.n609 2.2005
R15510 CLK_IN.n612 CLK_IN.n611 2.2005
R15511 CLK_IN.n514 CLK_IN.n513 2.2005
R15512 CLK_IN.n618 CLK_IN.n617 2.2005
R15513 CLK_IN.n620 CLK_IN.n512 2.2005
R15514 CLK_IN.n622 CLK_IN.n621 2.2005
R15515 CLK_IN.n625 CLK_IN.n624 2.2005
R15516 CLK_IN.n626 CLK_IN.n511 2.2005
R15517 CLK_IN.n628 CLK_IN.n627 2.2005
R15518 CLK_IN.n631 CLK_IN.n630 2.2005
R15519 CLK_IN.n629 CLK_IN.n509 2.2005
R15520 CLK_IN.n636 CLK_IN.n508 2.2005
R15521 CLK_IN.n639 CLK_IN.n638 2.2005
R15522 CLK_IN.n641 CLK_IN.n507 2.2005
R15523 CLK_IN.n643 CLK_IN.n642 2.2005
R15524 CLK_IN.n645 CLK_IN.n644 2.2005
R15525 CLK_IN.n498 CLK_IN.n496 2.2005
R15526 CLK_IN.n651 CLK_IN.n650 2.2005
R15527 CLK_IN.n505 CLK_IN.n497 2.2005
R15528 CLK_IN.n504 CLK_IN.n503 2.2005
R15529 CLK_IN.n502 CLK_IN.n501 2.2005
R15530 CLK_IN.n82 CLK_IN.n80 2.2005
R15531 CLK_IN.n1301 CLK_IN.n1300 2.2005
R15532 CLK_IN.n83 CLK_IN.n81 2.2005
R15533 CLK_IN.n823 CLK_IN.n822 2.2005
R15534 CLK_IN.n262 CLK_IN.n253 2.2005
R15535 CLK_IN.n263 CLK_IN.n257 2.2005
R15536 CLK_IN.n817 CLK_IN.n816 2.2005
R15537 CLK_IN.n260 CLK_IN.n258 2.2005
R15538 CLK_IN.n290 CLK_IN.n289 2.2005
R15539 CLK_IN.n292 CLK_IN.n291 2.2005
R15540 CLK_IN.n295 CLK_IN.n294 2.2005
R15541 CLK_IN.n296 CLK_IN.n272 2.2005
R15542 CLK_IN.n809 CLK_IN.n273 2.2005
R15543 CLK_IN.n807 CLK_IN.n806 2.2005
R15544 CLK_IN.n805 CLK_IN.n804 2.2005
R15545 CLK_IN.n802 CLK_IN.n801 2.2005
R15546 CLK_IN.n800 CLK_IN.n799 2.2005
R15547 CLK_IN.n797 CLK_IN.n796 2.2005
R15548 CLK_IN.n795 CLK_IN.n280 2.2005
R15549 CLK_IN.n311 CLK_IN.n281 2.2005
R15550 CLK_IN.n310 CLK_IN.n306 2.2005
R15551 CLK_IN.n790 CLK_IN.n789 2.2005
R15552 CLK_IN.n309 CLK_IN.n307 2.2005
R15553 CLK_IN.n323 CLK_IN.n322 2.2005
R15554 CLK_IN.n325 CLK_IN.n324 2.2005
R15555 CLK_IN.n319 CLK_IN.n317 2.2005
R15556 CLK_IN.n783 CLK_IN.n782 2.2005
R15557 CLK_IN.n320 CLK_IN.n318 2.2005
R15558 CLK_IN.n336 CLK_IN.n333 2.2005
R15559 CLK_IN.n777 CLK_IN.n776 2.2005
R15560 CLK_IN.n338 CLK_IN.n334 2.2005
R15561 CLK_IN.n771 CLK_IN.n342 2.2005
R15562 CLK_IN.n769 CLK_IN.n768 2.2005
R15563 CLK_IN.n352 CLK_IN.n344 2.2005
R15564 CLK_IN.n353 CLK_IN.n349 2.2005
R15565 CLK_IN.n763 CLK_IN.n762 2.2005
R15566 CLK_IN.n354 CLK_IN.n350 2.2005
R15567 CLK_IN.n360 CLK_IN.n358 2.2005
R15568 CLK_IN.n756 CLK_IN.n361 2.2005
R15569 CLK_IN.n754 CLK_IN.n753 2.2005
R15570 CLK_IN.n752 CLK_IN.n751 2.2005
R15571 CLK_IN.n750 CLK_IN.n749 2.2005
R15572 CLK_IN.n748 CLK_IN.n747 2.2005
R15573 CLK_IN.n745 CLK_IN.n744 2.2005
R15574 CLK_IN.n386 CLK_IN.n369 2.2005
R15575 CLK_IN.n387 CLK_IN.n380 2.2005
R15576 CLK_IN.n739 CLK_IN.n738 2.2005
R15577 CLK_IN.n383 CLK_IN.n381 2.2005
R15578 CLK_IN.n402 CLK_IN.n401 2.2005
R15579 CLK_IN.n404 CLK_IN.n403 2.2005
R15580 CLK_IN.n407 CLK_IN.n406 2.2005
R15581 CLK_IN.n405 CLK_IN.n394 2.2005
R15582 CLK_IN.n732 CLK_IN.n731 2.2005
R15583 CLK_IN.n730 CLK_IN.n395 2.2005
R15584 CLK_IN.n419 CLK_IN.n397 2.2005
R15585 CLK_IN.n421 CLK_IN.n415 2.2005
R15586 CLK_IN.n725 CLK_IN.n724 2.2005
R15587 CLK_IN.n423 CLK_IN.n416 2.2005
R15588 CLK_IN.n427 CLK_IN.n424 2.2005
R15589 CLK_IN.n719 CLK_IN.n718 2.2005
R15590 CLK_IN.n428 CLK_IN.n425 2.2005
R15591 CLK_IN.n437 CLK_IN.n433 2.2005
R15592 CLK_IN.n713 CLK_IN.n712 2.2005
R15593 CLK_IN.n436 CLK_IN.n434 2.2005
R15594 CLK_IN.n706 CLK_IN.n445 2.2005
R15595 CLK_IN.n705 CLK_IN.n704 2.2005
R15596 CLK_IN.n455 CLK_IN.n447 2.2005
R15597 CLK_IN.n456 CLK_IN.n452 2.2005
R15598 CLK_IN.n1137 CLK_IN.n1136 2.2005
R15599 CLK_IN.n1146 CLK_IN.n1145 2.2005
R15600 CLK_IN.n1148 CLK_IN.n1147 2.2005
R15601 CLK_IN.n1150 CLK_IN.n1149 2.2005
R15602 CLK_IN.n1152 CLK_IN.n1151 2.2005
R15603 CLK_IN.n1153 CLK_IN.n123 2.2005
R15604 CLK_IN.n1155 CLK_IN.n1154 2.2005
R15605 CLK_IN.n1158 CLK_IN.n1157 2.2005
R15606 CLK_IN.n1160 CLK_IN.n1159 2.2005
R15607 CLK_IN.n1162 CLK_IN.n1161 2.2005
R15608 CLK_IN.n1164 CLK_IN.n1163 2.2005
R15609 CLK_IN.n1166 CLK_IN.n1165 2.2005
R15610 CLK_IN.n1167 CLK_IN.n119 2.2005
R15611 CLK_IN.n1170 CLK_IN.n1169 2.2005
R15612 CLK_IN.n1172 CLK_IN.n118 2.2005
R15613 CLK_IN.n1174 CLK_IN.n1173 2.2005
R15614 CLK_IN.n1177 CLK_IN.n1176 2.2005
R15615 CLK_IN.n1175 CLK_IN.n116 2.2005
R15616 CLK_IN.n1185 CLK_IN.n1184 2.2005
R15617 CLK_IN.n1187 CLK_IN.n1186 2.2005
R15618 CLK_IN.n1189 CLK_IN.n1188 2.2005
R15619 CLK_IN.n1191 CLK_IN.n1190 2.2005
R15620 CLK_IN.n1193 CLK_IN.n1192 2.2005
R15621 CLK_IN.n1195 CLK_IN.n1194 2.2005
R15622 CLK_IN.n1197 CLK_IN.n1196 2.2005
R15623 CLK_IN.n1199 CLK_IN.n1198 2.2005
R15624 CLK_IN.n1201 CLK_IN.n1200 2.2005
R15625 CLK_IN.n1203 CLK_IN.n1202 2.2005
R15626 CLK_IN.n110 CLK_IN.n109 2.2005
R15627 CLK_IN.n1209 CLK_IN.n1208 2.2005
R15628 CLK_IN.n1211 CLK_IN.n108 2.2005
R15629 CLK_IN.n1213 CLK_IN.n1212 2.2005
R15630 CLK_IN.n1215 CLK_IN.n1214 2.2005
R15631 CLK_IN.n1217 CLK_IN.n1216 2.2005
R15632 CLK_IN.n1219 CLK_IN.n1218 2.2005
R15633 CLK_IN.n1221 CLK_IN.n1220 2.2005
R15634 CLK_IN.n106 CLK_IN.n105 2.2005
R15635 CLK_IN.n1227 CLK_IN.n1226 2.2005
R15636 CLK_IN.n1229 CLK_IN.n104 2.2005
R15637 CLK_IN.n1231 CLK_IN.n1230 2.2005
R15638 CLK_IN.n1234 CLK_IN.n1233 2.2005
R15639 CLK_IN.n1236 CLK_IN.n1235 2.2005
R15640 CLK_IN.n1238 CLK_IN.n1237 2.2005
R15641 CLK_IN.n102 CLK_IN.n101 2.2005
R15642 CLK_IN.n1244 CLK_IN.n1243 2.2005
R15643 CLK_IN.n1246 CLK_IN.n100 2.2005
R15644 CLK_IN.n1248 CLK_IN.n1247 2.2005
R15645 CLK_IN.n1251 CLK_IN.n1250 2.2005
R15646 CLK_IN.n1253 CLK_IN.n1252 2.2005
R15647 CLK_IN.n1256 CLK_IN.n1255 2.2005
R15648 CLK_IN.n1254 CLK_IN.n98 2.2005
R15649 CLK_IN.n1263 CLK_IN.n1262 2.2005
R15650 CLK_IN.n1265 CLK_IN.n1264 2.2005
R15651 CLK_IN.n1267 CLK_IN.n1266 2.2005
R15652 CLK_IN.n1269 CLK_IN.n1268 2.2005
R15653 CLK_IN.n1271 CLK_IN.n1270 2.2005
R15654 CLK_IN.n1273 CLK_IN.n1272 2.2005
R15655 CLK_IN.n1275 CLK_IN.n1274 2.2005
R15656 CLK_IN.n1277 CLK_IN.n1276 2.2005
R15657 CLK_IN.n93 CLK_IN.n92 2.2005
R15658 CLK_IN.n1283 CLK_IN.n1282 2.2005
R15659 CLK_IN.n1285 CLK_IN.n91 2.2005
R15660 CLK_IN.n1287 CLK_IN.n1286 2.2005
R15661 CLK_IN.n1290 CLK_IN.n1289 2.2005
R15662 CLK_IN.n1292 CLK_IN.n1291 2.2005
R15663 CLK_IN.n842 CLK_IN.n237 1.8005
R15664 CLK_IN.n239 CLK_IN.n238 1.8005
R15665 CLK_IN.n913 CLK_IN.n912 1.8005
R15666 CLK_IN.n918 CLK_IN.n917 1.8005
R15667 CLK_IN.n968 CLK_IN.n967 1.8005
R15668 CLK_IN.n973 CLK_IN.n972 1.8005
R15669 CLK_IN.n1381 CLK_IN.n14 1.8005
R15670 CLK_IN.n177 CLK_IN.n17 1.8005
R15671 CLK_IN.n1374 CLK_IN.n20 1.8005
R15672 CLK_IN.n163 CLK_IN.n22 1.8005
R15673 CLK_IN.n1368 CLK_IN.n25 1.8005
R15674 CLK_IN.n1095 CLK_IN.n27 1.8005
R15675 CLK_IN.n1362 CLK_IN.n30 1.8005
R15676 CLK_IN.n1303 CLK_IN.n1302 1.8005
R15677 CLK_IN.n653 CLK_IN.n652 1.8005
R15678 CLK_IN.n640 CLK_IN.n493 1.8005
R15679 CLK_IN.n659 CLK_IN.n491 1.8005
R15680 CLK_IN.n619 CLK_IN.n488 1.8005
R15681 CLK_IN.n665 CLK_IN.n486 1.8005
R15682 CLK_IN.n670 CLK_IN.n482 1.8005
R15683 CLK_IN.n672 CLK_IN.n480 1.8005
R15684 CLK_IN.n676 CLK_IN.n477 1.8005
R15685 CLK_IN.n678 CLK_IN.n475 1.8005
R15686 CLK_IN.n682 CLK_IN.n472 1.8005
R15687 CLK_IN.n684 CLK_IN.n470 1.8005
R15688 CLK_IN.n689 CLK_IN.n688 1.8005
R15689 CLK_IN.n1304 CLK_IN.n1303 1.8005
R15690 CLK_IN.n653 CLK_IN.n494 1.8005
R15691 CLK_IN.n656 CLK_IN.n493 1.8005
R15692 CLK_IN.n659 CLK_IN.n489 1.8005
R15693 CLK_IN.n662 CLK_IN.n488 1.8005
R15694 CLK_IN.n665 CLK_IN.n484 1.8005
R15695 CLK_IN.n670 CLK_IN.n669 1.8005
R15696 CLK_IN.n673 CLK_IN.n672 1.8005
R15697 CLK_IN.n676 CLK_IN.n675 1.8005
R15698 CLK_IN.n679 CLK_IN.n678 1.8005
R15699 CLK_IN.n682 CLK_IN.n681 1.8005
R15700 CLK_IN.n685 CLK_IN.n684 1.8005
R15701 CLK_IN.n688 CLK_IN.n687 1.8005
R15702 CLK_IN.n467 CLK_IN.n451 1.8005
R15703 CLK_IN.n699 CLK_IN.n451 1.8005
R15704 CLK_IN.n1307 CLK_IN.n77 1.8005
R15705 CLK_IN.n1307 CLK_IN.n1306 1.8005
R15706 CLK_IN.n869 CLK_IN.n237 1.8005
R15707 CLK_IN.n870 CLK_IN.n239 1.8005
R15708 CLK_IN.n914 CLK_IN.n913 1.8005
R15709 CLK_IN.n917 CLK_IN.n916 1.8005
R15710 CLK_IN.n969 CLK_IN.n968 1.8005
R15711 CLK_IN.n972 CLK_IN.n971 1.8005
R15712 CLK_IN.n1382 CLK_IN.n1381 1.8005
R15713 CLK_IN.n1377 CLK_IN.n17 1.8005
R15714 CLK_IN.n1374 CLK_IN.n18 1.8005
R15715 CLK_IN.n1371 CLK_IN.n22 1.8005
R15716 CLK_IN.n1368 CLK_IN.n23 1.8005
R15717 CLK_IN.n1365 CLK_IN.n27 1.8005
R15718 CLK_IN.n1362 CLK_IN.n28 1.8005
R15719 CLK_IN.n10 CLK_IN.n6 1.64317
R15720 CLK_IN.n241 CLK_IN.n240 1.5005
R15721 CLK_IN.n252 CLK_IN.n241 1.5005
R15722 CLK_IN.n1138 CLK_IN.n32 1.5005
R15723 CLK_IN.n1359 CLK_IN.n32 1.5005
R15724 CLK_IN.n1142 CLK_IN.n131 1.1125
R15725 CLK_IN.n711 CLK_IN.n710 1.10836
R15726 CLK_IN.n442 CLK_IN.n435 1.10443
R15727 CLK_IN.n696 CLK_IN.n457 1.10381
R15728 CLK_IN.n1141 CLK_IN.n132 1.10372
R15729 CLK_IN.n438 CLK_IN.n422 1.10339
R15730 CLK_IN.n706 CLK_IN.n443 1.10272
R15731 CLK_IN.n709 CLK_IN.n436 1.10272
R15732 CLK_IN.n441 CLK_IN.n437 1.10272
R15733 CLK_IN.n1145 CLK_IN.n1144 1.10263
R15734 CLK_IN.n1148 CLK_IN.n130 1.10263
R15735 CLK_IN.n1299 CLK_IN.n1298 1.1005
R15736 CLK_IN.n693 CLK_IN.n692 1.1005
R15737 CLK_IN.n535 CLK_IN.n458 1.1005
R15738 CLK_IN.n533 CLK_IN.n532 1.1005
R15739 CLK_IN.n531 CLK_IN.n530 1.1005
R15740 CLK_IN.n552 CLK_IN.n528 1.1005
R15741 CLK_IN.n561 CLK_IN.n560 1.1005
R15742 CLK_IN.n563 CLK_IN.n562 1.1005
R15743 CLK_IN.n569 CLK_IN.n525 1.1005
R15744 CLK_IN.n575 CLK_IN.n574 1.1005
R15745 CLK_IN.n577 CLK_IN.n576 1.1005
R15746 CLK_IN.n521 CLK_IN.n520 1.1005
R15747 CLK_IN.n594 CLK_IN.n593 1.1005
R15748 CLK_IN.n597 CLK_IN.n596 1.1005
R15749 CLK_IN.n595 CLK_IN.n517 1.1005
R15750 CLK_IN.n516 CLK_IN.n515 1.1005
R15751 CLK_IN.n614 CLK_IN.n613 1.1005
R15752 CLK_IN.n616 CLK_IN.n615 1.1005
R15753 CLK_IN.n623 CLK_IN.n510 1.1005
R15754 CLK_IN.n633 CLK_IN.n632 1.1005
R15755 CLK_IN.n635 CLK_IN.n634 1.1005
R15756 CLK_IN.n637 CLK_IN.n506 1.1005
R15757 CLK_IN.n647 CLK_IN.n646 1.1005
R15758 CLK_IN.n649 CLK_IN.n648 1.1005
R15759 CLK_IN.n499 CLK_IN.n84 1.1005
R15760 CLK_IN.n694 CLK_IN.n454 1.1005
R15761 CLK_IN.n264 CLK_IN.n261 1.1005
R15762 CLK_IN.n810 CLK_IN.n270 1.1005
R15763 CLK_IN.n772 CLK_IN.n339 1.1005
R15764 CLK_IN.n757 CLK_IN.n356 1.1005
R15765 CLK_IN.n388 CLK_IN.n385 1.1005
R15766 CLK_IN.n695 CLK_IN.n446 1.1005
R15767 CLK_IN.n708 CLK_IN.n707 1.1005
R15768 CLK_IN.n440 CLK_IN.n439 1.1005
R15769 CLK_IN.n721 CLK_IN.n720 1.1005
R15770 CLK_IN.n734 CLK_IN.n733 1.1005
R15771 CLK_IN.n390 CLK_IN.n389 1.1005
R15772 CLK_IN.n362 CLK_IN.n357 1.1005
R15773 CLK_IN.n759 CLK_IN.n758 1.1005
R15774 CLK_IN.n343 CLK_IN.n340 1.1005
R15775 CLK_IN.n774 CLK_IN.n773 1.1005
R15776 CLK_IN.n785 CLK_IN.n784 1.1005
R15777 CLK_IN.n313 CLK_IN.n312 1.1005
R15778 CLK_IN.n812 CLK_IN.n811 1.1005
R15779 CLK_IN.n815 CLK_IN.n814 1.1005
R15780 CLK_IN.n266 CLK_IN.n265 1.1005
R15781 CLK_IN.n826 CLK_IN.n825 1.1005
R15782 CLK_IN.n831 CLK_IN.n828 1.1005
R15783 CLK_IN.n824 CLK_IN.n250 1.1005
R15784 CLK_IN.n827 CLK_IN.n247 1.1005
R15785 CLK_IN.n1134 CLK_IN.n1133 1.1005
R15786 CLK_IN.n1125 CLK_IN.n1124 1.1005
R15787 CLK_IN.n1123 CLK_IN.n137 1.1005
R15788 CLK_IN.n1120 CLK_IN.n1119 1.1005
R15789 CLK_IN.n1116 CLK_IN.n1115 1.1005
R15790 CLK_IN.n1109 CLK_IN.n144 1.1005
R15791 CLK_IN.n1111 CLK_IN.n1110 1.1005
R15792 CLK_IN.n1108 CLK_IN.n143 1.1005
R15793 CLK_IN.n1103 CLK_IN.n1102 1.1005
R15794 CLK_IN.n1090 CLK_IN.n150 1.1005
R15795 CLK_IN.n1089 CLK_IN.n1088 1.1005
R15796 CLK_IN.n1087 CLK_IN.n151 1.1005
R15797 CLK_IN.n1082 CLK_IN.n153 1.1005
R15798 CLK_IN.n1081 CLK_IN.n1080 1.1005
R15799 CLK_IN.n1079 CLK_IN.n154 1.1005
R15800 CLK_IN.n1071 CLK_IN.n160 1.1005
R15801 CLK_IN.n1062 CLK_IN.n164 1.1005
R15802 CLK_IN.n1061 CLK_IN.n1060 1.1005
R15803 CLK_IN.n166 CLK_IN.n165 1.1005
R15804 CLK_IN.n1053 CLK_IN.n1052 1.1005
R15805 CLK_IN.n1051 CLK_IN.n169 1.1005
R15806 CLK_IN.n1050 CLK_IN.n1049 1.1005
R15807 CLK_IN.n1047 CLK_IN.n1046 1.1005
R15808 CLK_IN.n1042 CLK_IN.n171 1.1005
R15809 CLK_IN.n1039 CLK_IN.n172 1.1005
R15810 CLK_IN.n1036 CLK_IN.n173 1.1005
R15811 CLK_IN.n1030 CLK_IN.n174 1.1005
R15812 CLK_IN.n1029 CLK_IN.n1028 1.1005
R15813 CLK_IN.n176 CLK_IN.n175 1.1005
R15814 CLK_IN.n1021 CLK_IN.n1020 1.1005
R15815 CLK_IN.n1012 CLK_IN.n1011 1.1005
R15816 CLK_IN.n1010 CLK_IN.n182 1.1005
R15817 CLK_IN.n1007 CLK_IN.n1006 1.1005
R15818 CLK_IN.n1003 CLK_IN.n1002 1.1005
R15819 CLK_IN.n996 CLK_IN.n188 1.1005
R15820 CLK_IN.n998 CLK_IN.n997 1.1005
R15821 CLK_IN.n995 CLK_IN.n187 1.1005
R15822 CLK_IN.n987 CLK_IN.n193 1.1005
R15823 CLK_IN.n982 CLK_IN.n981 1.1005
R15824 CLK_IN.n980 CLK_IN.n195 1.1005
R15825 CLK_IN.n977 CLK_IN.n196 1.1005
R15826 CLK_IN.n951 CLK_IN.n950 1.1005
R15827 CLK_IN.n955 CLK_IN.n954 1.1005
R15828 CLK_IN.n956 CLK_IN.n947 1.1005
R15829 CLK_IN.n958 CLK_IN.n957 1.1005
R15830 CLK_IN.n963 CLK_IN.n205 1.1005
R15831 CLK_IN.n933 CLK_IN.n210 1.1005
R15832 CLK_IN.n935 CLK_IN.n934 1.1005
R15833 CLK_IN.n931 CLK_IN.n209 1.1005
R15834 CLK_IN.n926 CLK_IN.n925 1.1005
R15835 CLK_IN.n924 CLK_IN.n212 1.1005
R15836 CLK_IN.n923 CLK_IN.n922 1.1005
R15837 CLK_IN.n901 CLK_IN.n214 1.1005
R15838 CLK_IN.n903 CLK_IN.n902 1.1005
R15839 CLK_IN.n906 CLK_IN.n905 1.1005
R15840 CLK_IN.n909 CLK_IN.n908 1.1005
R15841 CLK_IN.n898 CLK_IN.n897 1.1005
R15842 CLK_IN.n896 CLK_IN.n225 1.1005
R15843 CLK_IN.n895 CLK_IN.n894 1.1005
R15844 CLK_IN.n228 CLK_IN.n227 1.1005
R15845 CLK_IN.n886 CLK_IN.n885 1.1005
R15846 CLK_IN.n884 CLK_IN.n230 1.1005
R15847 CLK_IN.n880 CLK_IN.n231 1.1005
R15848 CLK_IN.n879 CLK_IN.n878 1.1005
R15849 CLK_IN.n876 CLK_IN.n875 1.1005
R15850 CLK_IN.n847 CLK_IN.n846 1.1005
R15851 CLK_IN.n851 CLK_IN.n845 1.1005
R15852 CLK_IN.n853 CLK_IN.n852 1.1005
R15853 CLK_IN.n854 CLK_IN.n841 1.1005
R15854 CLK_IN.n859 CLK_IN.n839 1.1005
R15855 CLK_IN.n837 CLK_IN.n836 1.1005
R15856 CLK_IN.n835 CLK_IN.n246 1.1005
R15857 CLK_IN.n249 CLK_IN.n248 1.1005
R15858 CLK_IN.n829 CLK_IN.n249 1.1005
R15859 CLK_IN.n832 CLK_IN.n831 1.1005
R15860 CLK_IN.n834 CLK_IN.n833 1.1005
R15861 CLK_IN.n861 CLK_IN.n860 1.1005
R15862 CLK_IN.n862 CLK_IN.n245 1.1005
R15863 CLK_IN.n864 CLK_IN.n863 1.1005
R15864 CLK_IN.n838 CLK_IN.n244 1.1005
R15865 CLK_IN.n858 CLK_IN.n857 1.1005
R15866 CLK_IN.n856 CLK_IN.n855 1.1005
R15867 CLK_IN.n850 CLK_IN.n849 1.1005
R15868 CLK_IN.n235 CLK_IN.n234 1.1005
R15869 CLK_IN.n877 CLK_IN.n232 1.1005
R15870 CLK_IN.n883 CLK_IN.n882 1.1005
R15871 CLK_IN.n892 CLK_IN.n891 1.1005
R15872 CLK_IN.n893 CLK_IN.n226 1.1005
R15873 CLK_IN.n899 CLK_IN.n223 1.1005
R15874 CLK_IN.n907 CLK_IN.n224 1.1005
R15875 CLK_IN.n904 CLK_IN.n900 1.1005
R15876 CLK_IN.n921 CLK_IN.n213 1.1005
R15877 CLK_IN.n927 CLK_IN.n211 1.1005
R15878 CLK_IN.n930 CLK_IN.n929 1.1005
R15879 CLK_IN.n932 CLK_IN.n207 1.1005
R15880 CLK_IN.n965 CLK_IN.n964 1.1005
R15881 CLK_IN.n943 CLK_IN.n204 1.1005
R15882 CLK_IN.n942 CLK_IN.n941 1.1005
R15883 CLK_IN.n940 CLK_IN.n206 1.1005
R15884 CLK_IN.n962 CLK_IN.n961 1.1005
R15885 CLK_IN.n959 CLK_IN.n944 1.1005
R15886 CLK_IN.n953 CLK_IN.n948 1.1005
R15887 CLK_IN.n949 CLK_IN.n197 1.1005
R15888 CLK_IN.n979 CLK_IN.n978 1.1005
R15889 CLK_IN.n989 CLK_IN.n988 1.1005
R15890 CLK_IN.n986 CLK_IN.n192 1.1005
R15891 CLK_IN.n985 CLK_IN.n984 1.1005
R15892 CLK_IN.n983 CLK_IN.n194 1.1005
R15893 CLK_IN.n190 CLK_IN.n189 1.1005
R15894 CLK_IN.n994 CLK_IN.n993 1.1005
R15895 CLK_IN.n186 CLK_IN.n185 1.1005
R15896 CLK_IN.n1004 CLK_IN.n184 1.1005
R15897 CLK_IN.n1005 CLK_IN.n183 1.1005
R15898 CLK_IN.n1019 CLK_IN.n179 1.1005
R15899 CLK_IN.n1014 CLK_IN.n180 1.1005
R15900 CLK_IN.n1016 CLK_IN.n1015 1.1005
R15901 CLK_IN.n1013 CLK_IN.n181 1.1005
R15902 CLK_IN.n1022 CLK_IN.n178 1.1005
R15903 CLK_IN.n1024 CLK_IN.n1023 1.1005
R15904 CLK_IN.n1032 CLK_IN.n1031 1.1005
R15905 CLK_IN.n1038 CLK_IN.n1037 1.1005
R15906 CLK_IN.n1041 CLK_IN.n1040 1.1005
R15907 CLK_IN.n1048 CLK_IN.n170 1.1005
R15908 CLK_IN.n1054 CLK_IN.n168 1.1005
R15909 CLK_IN.n1056 CLK_IN.n1055 1.1005
R15910 CLK_IN.n1064 CLK_IN.n1063 1.1005
R15911 CLK_IN.n1073 CLK_IN.n1072 1.1005
R15912 CLK_IN.n1070 CLK_IN.n159 1.1005
R15913 CLK_IN.n1069 CLK_IN.n1068 1.1005
R15914 CLK_IN.n162 CLK_IN.n161 1.1005
R15915 CLK_IN.n158 CLK_IN.n157 1.1005
R15916 CLK_IN.n1078 CLK_IN.n1077 1.1005
R15917 CLK_IN.n1084 CLK_IN.n1083 1.1005
R15918 CLK_IN.n1086 CLK_IN.n1085 1.1005
R15919 CLK_IN.n1093 CLK_IN.n1092 1.1005
R15920 CLK_IN.n1101 CLK_IN.n146 1.1005
R15921 CLK_IN.n1100 CLK_IN.n1099 1.1005
R15922 CLK_IN.n1098 CLK_IN.n147 1.1005
R15923 CLK_IN.n1091 CLK_IN.n148 1.1005
R15924 CLK_IN.n1104 CLK_IN.n145 1.1005
R15925 CLK_IN.n1107 CLK_IN.n1106 1.1005
R15926 CLK_IN.n141 CLK_IN.n140 1.1005
R15927 CLK_IN.n1117 CLK_IN.n139 1.1005
R15928 CLK_IN.n1118 CLK_IN.n138 1.1005
R15929 CLK_IN.n1126 CLK_IN.n136 1.1005
R15930 CLK_IN.n1132 CLK_IN.n134 1.1005
R15931 CLK_IN.n135 CLK_IN.n133 1.1005
R15932 CLK_IN.n1129 CLK_IN.n1128 1.1005
R15933 CLK_IN.n86 CLK_IN.n85 1.1005
R15934 CLK_IN.n1296 CLK_IN.n1295 1.1005
R15935 CLK_IN.n1297 CLK_IN.n1296 1.1005
R15936 CLK_IN.n1131 CLK_IN.n135 1.1005
R15937 CLK_IN.n1130 CLK_IN.n1129 1.1005
R15938 CLK_IN.n1294 CLK_IN.n1293 1.1005
R15939 CLK_IN.n1288 CLK_IN.n87 1.1005
R15940 CLK_IN.n1281 CLK_IN.n1280 1.1005
R15941 CLK_IN.n1279 CLK_IN.n1278 1.1005
R15942 CLK_IN.n95 CLK_IN.n94 1.1005
R15943 CLK_IN.n1259 CLK_IN.n96 1.1005
R15944 CLK_IN.n1261 CLK_IN.n1260 1.1005
R15945 CLK_IN.n1258 CLK_IN.n1257 1.1005
R15946 CLK_IN.n1249 CLK_IN.n99 1.1005
R15947 CLK_IN.n1242 CLK_IN.n1241 1.1005
R15948 CLK_IN.n1240 CLK_IN.n1239 1.1005
R15949 CLK_IN.n1232 CLK_IN.n103 1.1005
R15950 CLK_IN.n1225 CLK_IN.n1224 1.1005
R15951 CLK_IN.n1223 CLK_IN.n1222 1.1005
R15952 CLK_IN.n1214 CLK_IN.n107 1.1005
R15953 CLK_IN.n1207 CLK_IN.n1206 1.1005
R15954 CLK_IN.n1205 CLK_IN.n1204 1.1005
R15955 CLK_IN.n112 CLK_IN.n111 1.1005
R15956 CLK_IN.n1180 CLK_IN.n113 1.1005
R15957 CLK_IN.n1181 CLK_IN.n115 1.1005
R15958 CLK_IN.n1183 CLK_IN.n1182 1.1005
R15959 CLK_IN.n1179 CLK_IN.n1178 1.1005
R15960 CLK_IN.n1168 CLK_IN.n117 1.1005
R15961 CLK_IN.n126 CLK_IN.n120 1.1005
R15962 CLK_IN.n127 CLK_IN.n121 1.1005
R15963 CLK_IN.n128 CLK_IN.n122 1.1005
R15964 CLK_IN.n129 CLK_IN.n124 1.1005
R15965 CLK_IN.n1143 CLK_IN.n125 1.1005
R15966 CLK_IN.n1140 CLK_IN.n1139 1.1005
R15967 CLK_IN.n1384 CLK_IN.n10 0.9025
R15968 CLK_IN.n252 CLK_IN.n247 0.733833
R15969 CLK_IN.n699 CLK_IN.n698 0.733833
R15970 CLK_IN.n1293 CLK_IN.n77 0.733833
R15971 CLK_IN.n1139 CLK_IN.n1138 0.733833
R15972 CLK_IN.n385 CLK_IN.n382 0.573769
R15973 CLK_IN.n808 CLK_IN.n270 0.573769
R15974 CLK_IN.n755 CLK_IN.n356 0.573695
R15975 CLK_IN.n261 CLK_IN.n259 0.573695
R15976 CLK_IN.n770 CLK_IN.n339 0.573346
R15977 CLK_IN.n831 CLK_IN.n830 0.550549
R15978 CLK_IN.n1127 CLK_IN.n135 0.550549
R15979 CLK_IN.n390 CLK_IN.n368 0.39244
R15980 CLK_IN.n812 CLK_IN.n269 0.39244
R15981 CLK_IN.n759 CLK_IN.n355 0.389994
R15982 CLK_IN.n266 CLK_IN.n251 0.389994
R15983 CLK_IN.n775 CLK_IN.n774 0.387191
R15984 CLK_IN.n723 CLK_IN.n722 0.384705
R15985 CLK_IN.n786 CLK_IN.n314 0.384705
R15986 CLK_IN.n736 CLK_IN.n384 0.384705
R15987 CLK_IN.n803 CLK_IN.n271 0.384705
R15988 CLK_IN.n420 CLK_IN.n393 0.382331
R15989 CLK_IN.n788 CLK_IN.n787 0.382331
R15990 CLK_IN.n735 CLK_IN.n391 0.382034
R15991 CLK_IN.n279 CLK_IN.n277 0.382034
R15992 CLK_IN.n367 CLK_IN.n365 0.379547
R15993 CLK_IN.n337 CLK_IN.n316 0.379547
R15994 CLK_IN.n813 CLK_IN.n267 0.379547
R15995 CLK_IN.n760 CLK_IN.n351 0.376968
R15996 CLK_IN.n761 CLK_IN.n760 0.376876
R15997 CLK_IN.n746 CLK_IN.n367 0.375976
R15998 CLK_IN.n813 CLK_IN.n268 0.375976
R15999 CLK_IN.n335 CLK_IN.n316 0.375884
R16000 CLK_IN.n735 CLK_IN.n392 0.374982
R16001 CLK_IN.n798 CLK_IN.n279 0.374982
R16002 CLK_IN.n418 CLK_IN.n393 0.374889
R16003 CLK_IN.n787 CLK_IN.n308 0.374889
R16004 CLK_IN.n722 CLK_IN.n417 0.373984
R16005 CLK_IN.n786 CLK_IN.n315 0.373984
R16006 CLK_IN.n737 CLK_IN.n736 0.373891
R16007 CLK_IN.n274 CLK_IN.n271 0.373891
R16008 CLK_IN.n698 CLK_IN.n697 0.275034
R16009 CLK_IN.n5 CLK_IN.n3 0.238833
R16010 CLK_IN CLK_IN.n1383 0.148744
R16011 CLK_IN CLK_IN.n1384 0.0489
R16012 CLK_IN.n867 CLK_IN.n237 0.0405
R16013 CLK_IN.n872 CLK_IN.n237 0.0405
R16014 CLK_IN.n872 CLK_IN.n239 0.0405
R16015 CLK_IN.n239 CLK_IN.n219 0.0405
R16016 CLK_IN.n913 CLK_IN.n219 0.0405
R16017 CLK_IN.n913 CLK_IN.n217 0.0405
R16018 CLK_IN.n917 CLK_IN.n217 0.0405
R16019 CLK_IN.n917 CLK_IN.n201 0.0405
R16020 CLK_IN.n968 CLK_IN.n201 0.0405
R16021 CLK_IN.n968 CLK_IN.n199 0.0405
R16022 CLK_IN.n972 CLK_IN.n199 0.0405
R16023 CLK_IN.n972 CLK_IN.n13 0.0405
R16024 CLK_IN.n1381 CLK_IN.n13 0.0405
R16025 CLK_IN.n1381 CLK_IN.n1380 0.0405
R16026 CLK_IN.n1379 CLK_IN.n17 0.0405
R16027 CLK_IN.n1375 CLK_IN.n17 0.0405
R16028 CLK_IN.n1375 CLK_IN.n1374 0.0405
R16029 CLK_IN.n1374 CLK_IN.n1373 0.0405
R16030 CLK_IN.n1373 CLK_IN.n22 0.0405
R16031 CLK_IN.n1369 CLK_IN.n22 0.0405
R16032 CLK_IN.n1369 CLK_IN.n1368 0.0405
R16033 CLK_IN.n1368 CLK_IN.n1367 0.0405
R16034 CLK_IN.n1367 CLK_IN.n27 0.0405
R16035 CLK_IN.n1363 CLK_IN.n27 0.0405
R16036 CLK_IN.n1363 CLK_IN.n1362 0.0405
R16037 CLK_IN.n1362 CLK_IN.n1361 0.0405
R16038 CLK_IN.n688 CLK_IN.n465 0.0405
R16039 CLK_IN.n688 CLK_IN.n466 0.0405
R16040 CLK_IN.n684 CLK_IN.n466 0.0405
R16041 CLK_IN.n684 CLK_IN.n683 0.0405
R16042 CLK_IN.n683 CLK_IN.n682 0.0405
R16043 CLK_IN.n682 CLK_IN.n473 0.0405
R16044 CLK_IN.n678 CLK_IN.n473 0.0405
R16045 CLK_IN.n678 CLK_IN.n677 0.0405
R16046 CLK_IN.n677 CLK_IN.n676 0.0405
R16047 CLK_IN.n676 CLK_IN.n478 0.0405
R16048 CLK_IN.n672 CLK_IN.n478 0.0405
R16049 CLK_IN.n672 CLK_IN.n671 0.0405
R16050 CLK_IN.n671 CLK_IN.n670 0.0405
R16051 CLK_IN.n670 CLK_IN.n483 0.0405
R16052 CLK_IN.n666 CLK_IN.n665 0.0405
R16053 CLK_IN.n665 CLK_IN.n664 0.0405
R16054 CLK_IN.n664 CLK_IN.n488 0.0405
R16055 CLK_IN.n660 CLK_IN.n488 0.0405
R16056 CLK_IN.n660 CLK_IN.n659 0.0405
R16057 CLK_IN.n659 CLK_IN.n658 0.0405
R16058 CLK_IN.n658 CLK_IN.n493 0.0405
R16059 CLK_IN.n654 CLK_IN.n493 0.0405
R16060 CLK_IN.n654 CLK_IN.n653 0.0405
R16061 CLK_IN.n653 CLK_IN.n79 0.0405
R16062 CLK_IN.n1303 CLK_IN.n79 0.0405
R16063 CLK_IN.n1303 CLK_IN.n76 0.0405
R16064 CLK_IN.n687 CLK_IN.n468 0.0405
R16065 CLK_IN.n687 CLK_IN.n686 0.0405
R16066 CLK_IN.n686 CLK_IN.n685 0.0405
R16067 CLK_IN.n685 CLK_IN.n469 0.0405
R16068 CLK_IN.n681 CLK_IN.n469 0.0405
R16069 CLK_IN.n681 CLK_IN.n680 0.0405
R16070 CLK_IN.n680 CLK_IN.n679 0.0405
R16071 CLK_IN.n679 CLK_IN.n474 0.0405
R16072 CLK_IN.n675 CLK_IN.n474 0.0405
R16073 CLK_IN.n675 CLK_IN.n674 0.0405
R16074 CLK_IN.n674 CLK_IN.n673 0.0405
R16075 CLK_IN.n673 CLK_IN.n479 0.0405
R16076 CLK_IN.n669 CLK_IN.n479 0.0405
R16077 CLK_IN.n669 CLK_IN.n668 0.0405
R16078 CLK_IN.n667 CLK_IN.n484 0.0405
R16079 CLK_IN.n663 CLK_IN.n484 0.0405
R16080 CLK_IN.n663 CLK_IN.n662 0.0405
R16081 CLK_IN.n662 CLK_IN.n661 0.0405
R16082 CLK_IN.n661 CLK_IN.n489 0.0405
R16083 CLK_IN.n657 CLK_IN.n489 0.0405
R16084 CLK_IN.n657 CLK_IN.n656 0.0405
R16085 CLK_IN.n656 CLK_IN.n655 0.0405
R16086 CLK_IN.n655 CLK_IN.n494 0.0405
R16087 CLK_IN.n494 CLK_IN.n78 0.0405
R16088 CLK_IN.n1304 CLK_IN.n78 0.0405
R16089 CLK_IN.n1305 CLK_IN.n1304 0.0405
R16090 CLK_IN.n869 CLK_IN.n868 0.0405
R16091 CLK_IN.n871 CLK_IN.n869 0.0405
R16092 CLK_IN.n871 CLK_IN.n870 0.0405
R16093 CLK_IN.n870 CLK_IN.n218 0.0405
R16094 CLK_IN.n914 CLK_IN.n218 0.0405
R16095 CLK_IN.n915 CLK_IN.n914 0.0405
R16096 CLK_IN.n916 CLK_IN.n915 0.0405
R16097 CLK_IN.n916 CLK_IN.n200 0.0405
R16098 CLK_IN.n969 CLK_IN.n200 0.0405
R16099 CLK_IN.n970 CLK_IN.n969 0.0405
R16100 CLK_IN.n971 CLK_IN.n970 0.0405
R16101 CLK_IN.n971 CLK_IN.n11 0.0405
R16102 CLK_IN.n1382 CLK_IN.n12 0.0405
R16103 CLK_IN.n1378 CLK_IN.n1377 0.0405
R16104 CLK_IN.n1377 CLK_IN.n1376 0.0405
R16105 CLK_IN.n1376 CLK_IN.n18 0.0405
R16106 CLK_IN.n1372 CLK_IN.n18 0.0405
R16107 CLK_IN.n1372 CLK_IN.n1371 0.0405
R16108 CLK_IN.n1371 CLK_IN.n1370 0.0405
R16109 CLK_IN.n1370 CLK_IN.n23 0.0405
R16110 CLK_IN.n1366 CLK_IN.n23 0.0405
R16111 CLK_IN.n1366 CLK_IN.n1365 0.0405
R16112 CLK_IN.n1365 CLK_IN.n1364 0.0405
R16113 CLK_IN.n1364 CLK_IN.n28 0.0405
R16114 CLK_IN.n1360 CLK_IN.n28 0.0405
R16115 CLK_IN.n1380 CLK_IN.n1379 0.0360676
R16116 CLK_IN.n666 CLK_IN.n483 0.0360676
R16117 CLK_IN.n668 CLK_IN.n667 0.0360676
R16118 CLK_IN.n255 CLK_IN.n254 0.0360676
R16119 CLK_IN.n285 CLK_IN.n255 0.0360676
R16120 CLK_IN.n286 CLK_IN.n285 0.0360676
R16121 CLK_IN.n287 CLK_IN.n286 0.0360676
R16122 CLK_IN.n287 CLK_IN.n283 0.0360676
R16123 CLK_IN.n301 CLK_IN.n283 0.0360676
R16124 CLK_IN.n302 CLK_IN.n301 0.0360676
R16125 CLK_IN.n303 CLK_IN.n302 0.0360676
R16126 CLK_IN.n304 CLK_IN.n303 0.0360676
R16127 CLK_IN.n328 CLK_IN.n304 0.0360676
R16128 CLK_IN.n329 CLK_IN.n328 0.0360676
R16129 CLK_IN.n330 CLK_IN.n329 0.0360676
R16130 CLK_IN.n331 CLK_IN.n330 0.0360676
R16131 CLK_IN.n345 CLK_IN.n331 0.0360676
R16132 CLK_IN.n346 CLK_IN.n345 0.0360676
R16133 CLK_IN.n347 CLK_IN.n346 0.0360676
R16134 CLK_IN.n371 CLK_IN.n347 0.0360676
R16135 CLK_IN.n372 CLK_IN.n371 0.0360676
R16136 CLK_IN.n375 CLK_IN.n372 0.0360676
R16137 CLK_IN.n376 CLK_IN.n375 0.0360676
R16138 CLK_IN.n377 CLK_IN.n376 0.0360676
R16139 CLK_IN.n378 CLK_IN.n377 0.0360676
R16140 CLK_IN.n399 CLK_IN.n378 0.0360676
R16141 CLK_IN.n410 CLK_IN.n399 0.0360676
R16142 CLK_IN.n411 CLK_IN.n410 0.0360676
R16143 CLK_IN.n412 CLK_IN.n411 0.0360676
R16144 CLK_IN.n413 CLK_IN.n412 0.0360676
R16145 CLK_IN.n429 CLK_IN.n413 0.0360676
R16146 CLK_IN.n430 CLK_IN.n429 0.0360676
R16147 CLK_IN.n431 CLK_IN.n430 0.0360676
R16148 CLK_IN.n448 CLK_IN.n431 0.0360676
R16149 CLK_IN.n449 CLK_IN.n448 0.0360676
R16150 CLK_IN.n450 CLK_IN.n449 0.0360676
R16151 CLK_IN.n820 CLK_IN.n819 0.0360676
R16152 CLK_IN.n819 CLK_IN.n256 0.0360676
R16153 CLK_IN.n284 CLK_IN.n256 0.0360676
R16154 CLK_IN.n298 CLK_IN.n284 0.0360676
R16155 CLK_IN.n299 CLK_IN.n298 0.0360676
R16156 CLK_IN.n300 CLK_IN.n299 0.0360676
R16157 CLK_IN.n300 CLK_IN.n282 0.0360676
R16158 CLK_IN.n793 CLK_IN.n282 0.0360676
R16159 CLK_IN.n793 CLK_IN.n792 0.0360676
R16160 CLK_IN.n792 CLK_IN.n305 0.0360676
R16161 CLK_IN.n327 CLK_IN.n305 0.0360676
R16162 CLK_IN.n780 CLK_IN.n327 0.0360676
R16163 CLK_IN.n780 CLK_IN.n779 0.0360676
R16164 CLK_IN.n779 CLK_IN.n332 0.0360676
R16165 CLK_IN.n766 CLK_IN.n332 0.0360676
R16166 CLK_IN.n766 CLK_IN.n765 0.0360676
R16167 CLK_IN.n765 CLK_IN.n348 0.0360676
R16168 CLK_IN.n373 CLK_IN.n348 0.0360676
R16169 CLK_IN.n374 CLK_IN.n373 0.0360676
R16170 CLK_IN.n374 CLK_IN.n370 0.0360676
R16171 CLK_IN.n742 CLK_IN.n370 0.0360676
R16172 CLK_IN.n742 CLK_IN.n741 0.0360676
R16173 CLK_IN.n741 CLK_IN.n379 0.0360676
R16174 CLK_IN.n409 CLK_IN.n379 0.0360676
R16175 CLK_IN.n409 CLK_IN.n398 0.0360676
R16176 CLK_IN.n728 CLK_IN.n398 0.0360676
R16177 CLK_IN.n728 CLK_IN.n727 0.0360676
R16178 CLK_IN.n727 CLK_IN.n414 0.0360676
R16179 CLK_IN.n716 CLK_IN.n414 0.0360676
R16180 CLK_IN.n716 CLK_IN.n715 0.0360676
R16181 CLK_IN.n715 CLK_IN.n432 0.0360676
R16182 CLK_IN.n702 CLK_IN.n432 0.0360676
R16183 CLK_IN.n702 CLK_IN.n701 0.0360676
R16184 CLK_IN.n1357 CLK_IN.n1356 0.0360676
R16185 CLK_IN.n1356 CLK_IN.n1355 0.0360676
R16186 CLK_IN.n1355 CLK_IN.n37 0.0360676
R16187 CLK_IN.n1351 CLK_IN.n37 0.0360676
R16188 CLK_IN.n1351 CLK_IN.n1350 0.0360676
R16189 CLK_IN.n1350 CLK_IN.n1349 0.0360676
R16190 CLK_IN.n1349 CLK_IN.n42 0.0360676
R16191 CLK_IN.n1345 CLK_IN.n42 0.0360676
R16192 CLK_IN.n1345 CLK_IN.n1344 0.0360676
R16193 CLK_IN.n1344 CLK_IN.n1343 0.0360676
R16194 CLK_IN.n1343 CLK_IN.n47 0.0360676
R16195 CLK_IN.n1339 CLK_IN.n47 0.0360676
R16196 CLK_IN.n1339 CLK_IN.n1338 0.0360676
R16197 CLK_IN.n1338 CLK_IN.n1337 0.0360676
R16198 CLK_IN.n1337 CLK_IN.n52 0.0360676
R16199 CLK_IN.n1333 CLK_IN.n52 0.0360676
R16200 CLK_IN.n1333 CLK_IN.n1332 0.0360676
R16201 CLK_IN.n1332 CLK_IN.n1331 0.0360676
R16202 CLK_IN.n1331 CLK_IN.n57 0.0360676
R16203 CLK_IN.n1327 CLK_IN.n57 0.0360676
R16204 CLK_IN.n1327 CLK_IN.n1326 0.0360676
R16205 CLK_IN.n1326 CLK_IN.n1325 0.0360676
R16206 CLK_IN.n1325 CLK_IN.n62 0.0360676
R16207 CLK_IN.n1321 CLK_IN.n62 0.0360676
R16208 CLK_IN.n1321 CLK_IN.n1320 0.0360676
R16209 CLK_IN.n1320 CLK_IN.n1319 0.0360676
R16210 CLK_IN.n1319 CLK_IN.n67 0.0360676
R16211 CLK_IN.n1315 CLK_IN.n67 0.0360676
R16212 CLK_IN.n1315 CLK_IN.n1314 0.0360676
R16213 CLK_IN.n1314 CLK_IN.n1313 0.0360676
R16214 CLK_IN.n1313 CLK_IN.n72 0.0360676
R16215 CLK_IN.n1309 CLK_IN.n72 0.0360676
R16216 CLK_IN.n1309 CLK_IN.n1308 0.0360676
R16217 CLK_IN.n1358 CLK_IN.n33 0.0360676
R16218 CLK_IN.n1354 CLK_IN.n33 0.0360676
R16219 CLK_IN.n1354 CLK_IN.n1353 0.0360676
R16220 CLK_IN.n1353 CLK_IN.n1352 0.0360676
R16221 CLK_IN.n1352 CLK_IN.n38 0.0360676
R16222 CLK_IN.n1348 CLK_IN.n38 0.0360676
R16223 CLK_IN.n1348 CLK_IN.n1347 0.0360676
R16224 CLK_IN.n1347 CLK_IN.n1346 0.0360676
R16225 CLK_IN.n1346 CLK_IN.n43 0.0360676
R16226 CLK_IN.n1342 CLK_IN.n43 0.0360676
R16227 CLK_IN.n1342 CLK_IN.n1341 0.0360676
R16228 CLK_IN.n1341 CLK_IN.n1340 0.0360676
R16229 CLK_IN.n1340 CLK_IN.n48 0.0360676
R16230 CLK_IN.n1336 CLK_IN.n48 0.0360676
R16231 CLK_IN.n1336 CLK_IN.n1335 0.0360676
R16232 CLK_IN.n1335 CLK_IN.n1334 0.0360676
R16233 CLK_IN.n1334 CLK_IN.n53 0.0360676
R16234 CLK_IN.n1330 CLK_IN.n53 0.0360676
R16235 CLK_IN.n1330 CLK_IN.n1329 0.0360676
R16236 CLK_IN.n1329 CLK_IN.n1328 0.0360676
R16237 CLK_IN.n1328 CLK_IN.n58 0.0360676
R16238 CLK_IN.n1324 CLK_IN.n58 0.0360676
R16239 CLK_IN.n1324 CLK_IN.n1323 0.0360676
R16240 CLK_IN.n1323 CLK_IN.n1322 0.0360676
R16241 CLK_IN.n1322 CLK_IN.n63 0.0360676
R16242 CLK_IN.n1318 CLK_IN.n63 0.0360676
R16243 CLK_IN.n1318 CLK_IN.n1317 0.0360676
R16244 CLK_IN.n1317 CLK_IN.n1316 0.0360676
R16245 CLK_IN.n1316 CLK_IN.n68 0.0360676
R16246 CLK_IN.n1312 CLK_IN.n68 0.0360676
R16247 CLK_IN.n1312 CLK_IN.n1311 0.0360676
R16248 CLK_IN.n1311 CLK_IN.n1310 0.0360676
R16249 CLK_IN.n1310 CLK_IN.n73 0.0360676
R16250 CLK_IN.n1378 CLK_IN.n12 0.0360676
R16251 CLK_IN.n1383 CLK_IN.n11 0.0281757
R16252 CLK_IN.n867 CLK_IN.n241 0.0234189
R16253 CLK_IN.n465 CLK_IN.n451 0.0234189
R16254 CLK_IN.n468 CLK_IN.n467 0.0234189
R16255 CLK_IN.n868 CLK_IN.n240 0.0234189
R16256 CLK_IN.n1361 CLK_IN.n32 0.0233108
R16257 CLK_IN.n1307 CLK_IN.n76 0.0233108
R16258 CLK_IN.n1306 CLK_IN.n1305 0.0233108
R16259 CLK_IN.n1360 CLK_IN.n1359 0.0233108
R16260 CLK_IN.n254 CLK_IN.n240 0.0227703
R16261 CLK_IN.n820 CLK_IN.n241 0.0227703
R16262 CLK_IN.n1357 CLK_IN.n32 0.0227703
R16263 CLK_IN.n1359 CLK_IN.n1358 0.0227703
R16264 CLK_IN.n844 CLK_IN.n236 0.0188784
R16265 CLK_IN.n874 CLK_IN.n233 0.0188784
R16266 CLK_IN.n887 CLK_IN.n229 0.0188784
R16267 CLK_IN.n889 CLK_IN.n220 0.0188784
R16268 CLK_IN.n911 CLK_IN.n222 0.0188784
R16269 CLK_IN.n936 CLK_IN.n208 0.0188784
R16270 CLK_IN.n938 CLK_IN.n202 0.0188784
R16271 CLK_IN.n966 CLK_IN.n203 0.0188784
R16272 CLK_IN.n946 CLK_IN.n198 0.0188784
R16273 CLK_IN.n976 CLK_IN.n975 0.0188784
R16274 CLK_IN.n990 CLK_IN.n191 0.0188784
R16275 CLK_IN.n1000 CLK_IN.n999 0.0188784
R16276 CLK_IN.n1009 CLK_IN.n1008 0.0188784
R16277 CLK_IN.n1018 CLK_IN.n1017 0.0188784
R16278 CLK_IN.n1027 CLK_IN.n1026 0.0188784
R16279 CLK_IN.n1034 CLK_IN.n1033 0.0188784
R16280 CLK_IN.n1044 CLK_IN.n1043 0.0188784
R16281 CLK_IN.n1058 CLK_IN.n167 0.0188784
R16282 CLK_IN.n1075 CLK_IN.n1074 0.0188784
R16283 CLK_IN.n156 CLK_IN.n155 0.0188784
R16284 CLK_IN.n1094 CLK_IN.n149 0.0188784
R16285 CLK_IN.n1097 CLK_IN.n1096 0.0188784
R16286 CLK_IN.n1112 CLK_IN.n142 0.0188784
R16287 CLK_IN.n538 CLK_IN.n537 0.0188784
R16288 CLK_IN.n542 CLK_IN.n541 0.0188784
R16289 CLK_IN.n546 CLK_IN.n545 0.0188784
R16290 CLK_IN.n550 CLK_IN.n549 0.0188784
R16291 CLK_IN.n555 CLK_IN.n554 0.0188784
R16292 CLK_IN.n567 CLK_IN.n566 0.0188784
R16293 CLK_IN.n572 CLK_IN.n571 0.0188784
R16294 CLK_IN.n579 CLK_IN.n523 0.0188784
R16295 CLK_IN.n582 CLK_IN.n581 0.0188784
R16296 CLK_IN.n586 CLK_IN.n585 0.0188784
R16297 CLK_IN.n591 CLK_IN.n589 0.0188784
R16298 CLK_IN.n599 CLK_IN.n598 0.0188784
R16299 CLK_IN.n603 CLK_IN.n602 0.0188784
R16300 CLK_IN.n607 CLK_IN.n606 0.0188784
R16301 CLK_IN.n611 CLK_IN.n610 0.0188784
R16302 CLK_IN.n618 CLK_IN.n513 0.0188784
R16303 CLK_IN.n621 CLK_IN.n620 0.0188784
R16304 CLK_IN.n626 CLK_IN.n625 0.0188784
R16305 CLK_IN.n639 CLK_IN.n508 0.0188784
R16306 CLK_IN.n642 CLK_IN.n641 0.0188784
R16307 CLK_IN.n644 CLK_IN.n496 0.0188784
R16308 CLK_IN.n651 CLK_IN.n497 0.0188784
R16309 CLK_IN.n503 CLK_IN.n502 0.0188784
R16310 CLK_IN.n822 CLK_IN.n252 0.0188784
R16311 CLK_IN.n257 CLK_IN.n253 0.0188784
R16312 CLK_IN.n817 CLK_IN.n258 0.0188784
R16313 CLK_IN.n292 CLK_IN.n290 0.0188784
R16314 CLK_IN.n763 CLK_IN.n350 0.0188784
R16315 CLK_IN.n361 CLK_IN.n360 0.0188784
R16316 CLK_IN.n753 CLK_IN.n752 0.0188784
R16317 CLK_IN.n749 CLK_IN.n748 0.0188784
R16318 CLK_IN.n1138 CLK_IN.n1137 0.0188784
R16319 CLK_IN.n1147 CLK_IN.n1146 0.0188784
R16320 CLK_IN.n1151 CLK_IN.n1150 0.0188784
R16321 CLK_IN.n1155 CLK_IN.n123 0.0188784
R16322 CLK_IN.n1216 CLK_IN.n1215 0.0188784
R16323 CLK_IN.n1220 CLK_IN.n1219 0.0188784
R16324 CLK_IN.n1227 CLK_IN.n105 0.0188784
R16325 CLK_IN.n1230 CLK_IN.n1229 0.0188784
R16326 CLK_IN.n865 CLK_IN.n243 0.0187703
R16327 CLK_IN.n844 CLK_IN.n843 0.0187703
R16328 CLK_IN.n919 CLK_IN.n215 0.0187703
R16329 CLK_IN.n216 CLK_IN.n208 0.0187703
R16330 CLK_IN.n991 CLK_IN.n990 0.0187703
R16331 CLK_IN.n1059 CLK_IN.n1058 0.0187703
R16332 CLK_IN.n1067 CLK_IN.n1066 0.0187703
R16333 CLK_IN.n1113 CLK_IN.n1112 0.0187703
R16334 CLK_IN.n1122 CLK_IN.n1121 0.0187703
R16335 CLK_IN.n690 CLK_IN.n462 0.0187703
R16336 CLK_IN.n537 CLK_IN.n463 0.0187703
R16337 CLK_IN.n558 CLK_IN.n557 0.0187703
R16338 CLK_IN.n566 CLK_IN.n565 0.0187703
R16339 CLK_IN.n591 CLK_IN.n590 0.0187703
R16340 CLK_IN.n627 CLK_IN.n626 0.0187703
R16341 CLK_IN.n630 CLK_IN.n629 0.0187703
R16342 CLK_IN.n502 CLK_IN.n80 0.0187703
R16343 CLK_IN.n1301 CLK_IN.n81 0.0187703
R16344 CLK_IN.n296 CLK_IN.n273 0.0187703
R16345 CLK_IN.n806 CLK_IN.n805 0.0187703
R16346 CLK_IN.n801 CLK_IN.n800 0.0187703
R16347 CLK_IN.n796 CLK_IN.n795 0.0187703
R16348 CLK_IN.n306 CLK_IN.n281 0.0187703
R16349 CLK_IN.n790 CLK_IN.n307 0.0187703
R16350 CLK_IN.n325 CLK_IN.n323 0.0187703
R16351 CLK_IN.n782 CLK_IN.n319 0.0187703
R16352 CLK_IN.n333 CLK_IN.n320 0.0187703
R16353 CLK_IN.n777 CLK_IN.n334 0.0187703
R16354 CLK_IN.n768 CLK_IN.n342 0.0187703
R16355 CLK_IN.n349 CLK_IN.n344 0.0187703
R16356 CLK_IN.n380 CLK_IN.n369 0.0187703
R16357 CLK_IN.n739 CLK_IN.n381 0.0187703
R16358 CLK_IN.n404 CLK_IN.n402 0.0187703
R16359 CLK_IN.n407 CLK_IN.n405 0.0187703
R16360 CLK_IN.n731 CLK_IN.n730 0.0187703
R16361 CLK_IN.n415 CLK_IN.n397 0.0187703
R16362 CLK_IN.n725 CLK_IN.n416 0.0187703
R16363 CLK_IN.n718 CLK_IN.n427 0.0187703
R16364 CLK_IN.n433 CLK_IN.n428 0.0187703
R16365 CLK_IN.n713 CLK_IN.n434 0.0187703
R16366 CLK_IN.n704 CLK_IN.n445 0.0187703
R16367 CLK_IN.n452 CLK_IN.n447 0.0187703
R16368 CLK_IN.n1161 CLK_IN.n1160 0.0187703
R16369 CLK_IN.n1165 CLK_IN.n1164 0.0187703
R16370 CLK_IN.n1170 CLK_IN.n119 0.0187703
R16371 CLK_IN.n1173 CLK_IN.n1172 0.0187703
R16372 CLK_IN.n1176 CLK_IN.n1175 0.0187703
R16373 CLK_IN.n1186 CLK_IN.n1185 0.0187703
R16374 CLK_IN.n1190 CLK_IN.n1189 0.0187703
R16375 CLK_IN.n1194 CLK_IN.n1193 0.0187703
R16376 CLK_IN.n1198 CLK_IN.n1197 0.0187703
R16377 CLK_IN.n1202 CLK_IN.n1201 0.0187703
R16378 CLK_IN.n1209 CLK_IN.n109 0.0187703
R16379 CLK_IN.n1212 CLK_IN.n1211 0.0187703
R16380 CLK_IN.n1237 CLK_IN.n1236 0.0187703
R16381 CLK_IN.n1244 CLK_IN.n101 0.0187703
R16382 CLK_IN.n1247 CLK_IN.n1246 0.0187703
R16383 CLK_IN.n1252 CLK_IN.n1251 0.0187703
R16384 CLK_IN.n1255 CLK_IN.n1254 0.0187703
R16385 CLK_IN.n1264 CLK_IN.n1263 0.0187703
R16386 CLK_IN.n1268 CLK_IN.n1267 0.0187703
R16387 CLK_IN.n1272 CLK_IN.n1271 0.0187703
R16388 CLK_IN.n1276 CLK_IN.n1275 0.0187703
R16389 CLK_IN.n1283 CLK_IN.n92 0.0187703
R16390 CLK_IN.n1286 CLK_IN.n1285 0.0187703
R16391 CLK_IN.n1291 CLK_IN.n1290 0.0187703
R16392 CLK_IN.n874 CLK_IN.n873 0.0185541
R16393 CLK_IN.n1096 CLK_IN.n29 0.0185541
R16394 CLK_IN.n541 CLK_IN.n534 0.0185541
R16395 CLK_IN.n500 CLK_IN.n497 0.0185541
R16396 CLK_IN.n297 CLK_IN.n295 0.0184459
R16397 CLK_IN.n744 CLK_IN.n743 0.0184459
R16398 CLK_IN.n1157 CLK_IN.n39 0.0184459
R16399 CLK_IN.n1233 CLK_IN.n60 0.0184459
R16400 CLK_IN.n999 CLK_IN.n14 0.0182297
R16401 CLK_IN.n598 CLK_IN.n482 0.0182297
R16402 CLK_IN.n295 CLK_IN.n293 0.0181216
R16403 CLK_IN.n744 CLK_IN.n366 0.0181216
R16404 CLK_IN.n1157 CLK_IN.n1156 0.0181216
R16405 CLK_IN.n1233 CLK_IN.n59 0.0181216
R16406 CLK_IN.n919 CLK_IN.n918 0.0175811
R16407 CLK_IN.n1066 CLK_IN.n163 0.0175811
R16408 CLK_IN.n557 CLK_IN.n475 0.0175811
R16409 CLK_IN.n630 CLK_IN.n491 0.0175811
R16410 CLK_IN.n275 CLK_IN.n273 0.0173649
R16411 CLK_IN.n740 CLK_IN.n380 0.0173649
R16412 CLK_IN.n1161 CLK_IN.n40 0.0173649
R16413 CLK_IN.n1237 CLK_IN.n61 0.0173649
R16414 CLK_IN.n290 CLK_IN.n288 0.0170405
R16415 CLK_IN.n749 CLK_IN.n364 0.0170405
R16416 CLK_IN.n123 CLK_IN.n36 0.0170405
R16417 CLK_IN.n1229 CLK_IN.n1228 0.0170405
R16418 CLK_IN.n938 CLK_IN.n937 0.0167162
R16419 CLK_IN.n1044 CLK_IN.n21 0.0167162
R16420 CLK_IN.n571 CLK_IN.n476 0.0167162
R16421 CLK_IN.n621 CLK_IN.n490 0.0167162
R16422 CLK_IN.n805 CLK_IN.n276 0.0162838
R16423 CLK_IN.n400 CLK_IN.n381 0.0162838
R16424 CLK_IN.n1165 CLK_IN.n41 0.0162838
R16425 CLK_IN.n1245 CLK_IN.n1244 0.0162838
R16426 CLK_IN.n975 CLK_IN.n974 0.0159595
R16427 CLK_IN.n1017 CLK_IN.n16 0.0159595
R16428 CLK_IN.n586 CLK_IN.n481 0.0159595
R16429 CLK_IN.n606 CLK_IN.n485 0.0159595
R16430 CLK_IN.n818 CLK_IN.n817 0.0159595
R16431 CLK_IN.n753 CLK_IN.n363 0.0159595
R16432 CLK_IN.n1150 CLK_IN.n35 0.0159595
R16433 CLK_IN.n105 CLK_IN.n56 0.0159595
R16434 CLK_IN.n842 CLK_IN.n243 0.0157432
R16435 CLK_IN.n1121 CLK_IN.n30 0.0157432
R16436 CLK_IN.n690 CLK_IN.n689 0.0157432
R16437 CLK_IN.n1302 CLK_IN.n1301 0.0157432
R16438 CLK_IN.n238 CLK_IN.n229 0.0152027
R16439 CLK_IN.n1095 CLK_IN.n1094 0.0152027
R16440 CLK_IN.n545 CLK_IN.n470 0.0152027
R16441 CLK_IN.n652 CLK_IN.n496 0.0152027
R16442 CLK_IN.n800 CLK_IN.n278 0.0152027
R16443 CLK_IN.n408 CLK_IN.n404 0.0152027
R16444 CLK_IN.n1171 CLK_IN.n1170 0.0152027
R16445 CLK_IN.n1247 CLK_IN.n64 0.0152027
R16446 CLK_IN.n1008 CLK_IN.n15 0.0148784
R16447 CLK_IN.n602 CLK_IN.n518 0.0148784
R16448 CLK_IN.n821 CLK_IN.n253 0.0148784
R16449 CLK_IN.n360 CLK_IN.n359 0.0148784
R16450 CLK_IN.n1146 CLK_IN.n34 0.0148784
R16451 CLK_IN.n1219 CLK_IN.n55 0.0148784
R16452 CLK_IN.n222 CLK_IN.n221 0.0141216
R16453 CLK_IN.n1074 CLK_IN.n24 0.0141216
R16454 CLK_IN.n556 CLK_IN.n555 0.0141216
R16455 CLK_IN.n508 CLK_IN.n492 0.0141216
R16456 CLK_IN.n795 CLK_IN.n794 0.0141216
R16457 CLK_IN.n405 CLK_IN.n396 0.0141216
R16458 CLK_IN.n1173 CLK_IN.n44 0.0141216
R16459 CLK_IN.n1252 CLK_IN.n65 0.0141216
R16460 CLK_IN.n467 CLK_IN.n450 0.0137973
R16461 CLK_IN.n701 CLK_IN.n451 0.0137973
R16462 CLK_IN.n764 CLK_IN.n763 0.0137973
R16463 CLK_IN.n700 CLK_IN.n699 0.0137973
R16464 CLK_IN.n1215 CLK_IN.n54 0.0137973
R16465 CLK_IN.n77 CLK_IN.n75 0.0137973
R16466 CLK_IN.n1308 CLK_IN.n1307 0.0137973
R16467 CLK_IN.n1306 CLK_IN.n73 0.0137973
R16468 CLK_IN.n1294 CLK_IN.n87 0.0134381
R16469 CLK_IN.n967 CLK_IN.n966 0.0133649
R16470 CLK_IN.n1033 CLK_IN.n20 0.0133649
R16471 CLK_IN.n523 CLK_IN.n477 0.0133649
R16472 CLK_IN.n619 CLK_IN.n618 0.0133649
R16473 CLK_IN.n791 CLK_IN.n306 0.0130405
R16474 CLK_IN.n730 CLK_IN.n729 0.0130405
R16475 CLK_IN.n1175 CLK_IN.n45 0.0130405
R16476 CLK_IN.n1254 CLK_IN.n66 0.0130405
R16477 CLK_IN.n767 CLK_IN.n344 0.0128243
R16478 CLK_IN.n703 CLK_IN.n447 0.0128243
R16479 CLK_IN.n1211 CLK_IN.n1210 0.0128243
R16480 CLK_IN.n1290 CLK_IN.n74 0.0128243
R16481 CLK_IN.n1383 CLK_IN.n1382 0.0128243
R16482 CLK_IN.n973 CLK_IN.n198 0.0126081
R16483 CLK_IN.n1026 CLK_IN.n177 0.0126081
R16484 CLK_IN.n582 CLK_IN.n480 0.0126081
R16485 CLK_IN.n610 CLK_IN.n486 0.0126081
R16486 CLK_IN.n866 CLK_IN.n242 0.0123919
R16487 CLK_IN.n1135 CLK_IN.n31 0.0123919
R16488 CLK_IN.n464 CLK_IN.n453 0.0123919
R16489 CLK_IN.n89 CLK_IN.n88 0.0123919
R16490 CLK_IN.n321 CLK_IN.n307 0.0119595
R16491 CLK_IN.n726 CLK_IN.n415 0.0119595
R16492 CLK_IN.n1186 CLK_IN.n46 0.0119595
R16493 CLK_IN.n1264 CLK_IN.n97 0.0119595
R16494 CLK_IN.n889 CLK_IN.n888 0.0118514
R16495 CLK_IN.n155 CLK_IN.n26 0.0118514
R16496 CLK_IN.n549 CLK_IN.n471 0.0118514
R16497 CLK_IN.n642 CLK_IN.n495 0.0118514
R16498 CLK_IN.n342 CLK_IN.n341 0.0117432
R16499 CLK_IN.n445 CLK_IN.n444 0.0117432
R16500 CLK_IN.n109 CLK_IN.n51 0.0117432
R16501 CLK_IN.n1285 CLK_IN.n1284 0.0117432
R16502 CLK_IN.n697 CLK_IN.n694 0.0116588
R16503 CLK_IN.n252 CLK_IN.n242 0.011527
R16504 CLK_IN.n699 CLK_IN.n453 0.011527
R16505 CLK_IN.n1138 CLK_IN.n1135 0.0114189
R16506 CLK_IN.n89 CLK_IN.n77 0.0114189
R16507 CLK_IN.n129 CLK_IN.n128 0.0109762
R16508 CLK_IN.n127 CLK_IN.n126 0.0109762
R16509 CLK_IN.n1179 CLK_IN.n117 0.0109762
R16510 CLK_IN.n1182 CLK_IN.n1181 0.0109762
R16511 CLK_IN.n1180 CLK_IN.n111 0.0109762
R16512 CLK_IN.n1206 CLK_IN.n1205 0.0109762
R16513 CLK_IN.n1223 CLK_IN.n107 0.0109762
R16514 CLK_IN.n1224 CLK_IN.n103 0.0109762
R16515 CLK_IN.n1241 CLK_IN.n1240 0.0109762
R16516 CLK_IN.n1258 CLK_IN.n99 0.0109762
R16517 CLK_IN.n1260 CLK_IN.n1259 0.0109762
R16518 CLK_IN.n1279 CLK_IN.n94 0.0109762
R16519 CLK_IN.n1280 CLK_IN.n87 0.0109762
R16520 CLK_IN.n693 CLK_IN.n458 0.0109762
R16521 CLK_IN.n532 CLK_IN.n458 0.0109762
R16522 CLK_IN.n532 CLK_IN.n531 0.0109762
R16523 CLK_IN.n531 CLK_IN.n528 0.0109762
R16524 CLK_IN.n561 CLK_IN.n528 0.0109762
R16525 CLK_IN.n562 CLK_IN.n561 0.0109762
R16526 CLK_IN.n562 CLK_IN.n525 0.0109762
R16527 CLK_IN.n575 CLK_IN.n525 0.0109762
R16528 CLK_IN.n576 CLK_IN.n575 0.0109762
R16529 CLK_IN.n576 CLK_IN.n520 0.0109762
R16530 CLK_IN.n594 CLK_IN.n520 0.0109762
R16531 CLK_IN.n596 CLK_IN.n595 0.0109762
R16532 CLK_IN.n595 CLK_IN.n515 0.0109762
R16533 CLK_IN.n614 CLK_IN.n515 0.0109762
R16534 CLK_IN.n615 CLK_IN.n614 0.0109762
R16535 CLK_IN.n615 CLK_IN.n510 0.0109762
R16536 CLK_IN.n633 CLK_IN.n510 0.0109762
R16537 CLK_IN.n634 CLK_IN.n633 0.0109762
R16538 CLK_IN.n634 CLK_IN.n506 0.0109762
R16539 CLK_IN.n647 CLK_IN.n506 0.0109762
R16540 CLK_IN.n648 CLK_IN.n647 0.0109762
R16541 CLK_IN.n648 CLK_IN.n84 0.0109762
R16542 CLK_IN.n1298 CLK_IN.n84 0.0109762
R16543 CLK_IN.n814 CLK_IN.n813 0.0109762
R16544 CLK_IN.n812 CLK_IN.n271 0.0109762
R16545 CLK_IN.n313 CLK_IN.n279 0.0109762
R16546 CLK_IN.n787 CLK_IN.n786 0.0109762
R16547 CLK_IN.n785 CLK_IN.n316 0.0109762
R16548 CLK_IN.n774 CLK_IN.n340 0.0109762
R16549 CLK_IN.n760 CLK_IN.n759 0.0109762
R16550 CLK_IN.n367 CLK_IN.n357 0.0109762
R16551 CLK_IN.n736 CLK_IN.n390 0.0109762
R16552 CLK_IN.n735 CLK_IN.n734 0.0109762
R16553 CLK_IN.n722 CLK_IN.n393 0.0109762
R16554 CLK_IN.n128 CLK_IN.n127 0.01095
R16555 CLK_IN.n126 CLK_IN.n117 0.01095
R16556 CLK_IN.n1182 CLK_IN.n1179 0.01095
R16557 CLK_IN.n1181 CLK_IN.n1180 0.01095
R16558 CLK_IN.n1205 CLK_IN.n111 0.01095
R16559 CLK_IN.n1206 CLK_IN.n107 0.01095
R16560 CLK_IN.n1224 CLK_IN.n1223 0.01095
R16561 CLK_IN.n1240 CLK_IN.n103 0.01095
R16562 CLK_IN.n1241 CLK_IN.n99 0.01095
R16563 CLK_IN.n1260 CLK_IN.n1258 0.01095
R16564 CLK_IN.n1259 CLK_IN.n94 0.01095
R16565 CLK_IN.n1280 CLK_IN.n1279 0.01095
R16566 CLK_IN.n596 CLK_IN.n594 0.01095
R16567 CLK_IN.n1298 CLK_IN.n1297 0.01095
R16568 CLK_IN.n814 CLK_IN.n266 0.01095
R16569 CLK_IN.n813 CLK_IN.n812 0.01095
R16570 CLK_IN.n279 CLK_IN.n271 0.01095
R16571 CLK_IN.n787 CLK_IN.n313 0.01095
R16572 CLK_IN.n786 CLK_IN.n785 0.01095
R16573 CLK_IN.n774 CLK_IN.n316 0.01095
R16574 CLK_IN.n760 CLK_IN.n340 0.01095
R16575 CLK_IN.n759 CLK_IN.n357 0.01095
R16576 CLK_IN.n390 CLK_IN.n367 0.01095
R16577 CLK_IN.n736 CLK_IN.n735 0.01095
R16578 CLK_IN.n734 CLK_IN.n393 0.01095
R16579 CLK_IN.n722 CLK_IN.n721 0.01095
R16580 CLK_IN.n326 CLK_IN.n325 0.0108784
R16581 CLK_IN.n426 CLK_IN.n416 0.0108784
R16582 CLK_IN.n1190 CLK_IN.n114 0.0108784
R16583 CLK_IN.n1268 CLK_IN.n69 0.0108784
R16584 CLK_IN.n912 CLK_IN.n220 0.0107703
R16585 CLK_IN.n156 CLK_IN.n25 0.0107703
R16586 CLK_IN.n550 CLK_IN.n472 0.0107703
R16587 CLK_IN.n641 CLK_IN.n640 0.0107703
R16588 CLK_IN.n778 CLK_IN.n777 0.0106622
R16589 CLK_IN.n714 CLK_IN.n713 0.0106622
R16590 CLK_IN.n1201 CLK_IN.n50 0.0106622
R16591 CLK_IN.n92 CLK_IN.n71 0.0106622
R16592 CLK_IN.n694 CLK_IN.n693 0.0106095
R16593 CLK_IN.n946 CLK_IN.n945 0.0100135
R16594 CLK_IN.n1027 CLK_IN.n19 0.0100135
R16595 CLK_IN.n581 CLK_IN.n580 0.0100135
R16596 CLK_IN.n611 CLK_IN.n487 0.0100135
R16597 CLK_IN.n782 CLK_IN.n781 0.0097973
R16598 CLK_IN.n718 CLK_IN.n717 0.0097973
R16599 CLK_IN.n1194 CLK_IN.n49 0.0097973
R16600 CLK_IN.n1272 CLK_IN.n70 0.0097973
R16601 CLK_IN.n697 CLK_IN.n696 0.00967266
R16602 CLK_IN.n781 CLK_IN.n320 0.00958108
R16603 CLK_IN.n717 CLK_IN.n428 0.00958108
R16604 CLK_IN.n1197 CLK_IN.n49 0.00958108
R16605 CLK_IN.n1275 CLK_IN.n70 0.00958108
R16606 CLK_IN.n945 CLK_IN.n203 0.00925676
R16607 CLK_IN.n1034 CLK_IN.n19 0.00925676
R16608 CLK_IN.n580 CLK_IN.n579 0.00925676
R16609 CLK_IN.n513 CLK_IN.n487 0.00925676
R16610 CLK_IN.n774 CLK_IN.n339 0.00880612
R16611 CLK_IN.n778 CLK_IN.n333 0.00871622
R16612 CLK_IN.n714 CLK_IN.n433 0.00871622
R16613 CLK_IN.n1198 CLK_IN.n50 0.00871622
R16614 CLK_IN.n1276 CLK_IN.n71 0.00871622
R16615 CLK_IN.n912 CLK_IN.n911 0.0085
R16616 CLK_IN.n1075 CLK_IN.n25 0.0085
R16617 CLK_IN.n554 CLK_IN.n472 0.0085
R16618 CLK_IN.n640 CLK_IN.n639 0.0085
R16619 CLK_IN.n326 CLK_IN.n319 0.0085
R16620 CLK_IN.n427 CLK_IN.n426 0.0085
R16621 CLK_IN.n1193 CLK_IN.n114 0.0085
R16622 CLK_IN.n1271 CLK_IN.n69 0.0085
R16623 CLK_IN.n130 CLK_IN.n129 0.00809524
R16624 CLK_IN.n695 CLK_IN.n443 0.00778095
R16625 CLK_IN.n341 CLK_IN.n334 0.00763514
R16626 CLK_IN.n444 CLK_IN.n434 0.00763514
R16627 CLK_IN.n1202 CLK_IN.n51 0.00763514
R16628 CLK_IN.n1284 CLK_IN.n1283 0.00763514
R16629 CLK_IN.n888 CLK_IN.n887 0.00741892
R16630 CLK_IN.n149 CLK_IN.n26 0.00741892
R16631 CLK_IN.n546 CLK_IN.n471 0.00741892
R16632 CLK_IN.n644 CLK_IN.n495 0.00741892
R16633 CLK_IN.n323 CLK_IN.n321 0.00741892
R16634 CLK_IN.n726 CLK_IN.n725 0.00741892
R16635 CLK_IN.n1189 CLK_IN.n46 0.00741892
R16636 CLK_IN.n1267 CLK_IN.n97 0.00741892
R16637 CLK_IN.n721 CLK_IN.n422 0.00725714
R16638 CLK_IN.n696 CLK_IN.n695 0.00707381
R16639 CLK_IN.n866 CLK_IN.n865 0.00698649
R16640 CLK_IN.n1122 CLK_IN.n31 0.00698649
R16641 CLK_IN.n464 CLK_IN.n462 0.00698649
R16642 CLK_IN.n88 CLK_IN.n81 0.00698649
R16643 CLK_IN.n266 CLK_IN.n250 0.00696162
R16644 CLK_IN.n1297 CLK_IN.n85 0.00691667
R16645 CLK_IN.n976 CLK_IN.n973 0.00666216
R16646 CLK_IN.n1018 CLK_IN.n177 0.00666216
R16647 CLK_IN.n585 CLK_IN.n480 0.00666216
R16648 CLK_IN.n607 CLK_IN.n486 0.00666216
R16649 CLK_IN.n768 CLK_IN.n767 0.00655405
R16650 CLK_IN.n704 CLK_IN.n703 0.00655405
R16651 CLK_IN.n1210 CLK_IN.n1209 0.00655405
R16652 CLK_IN.n1286 CLK_IN.n74 0.00655405
R16653 CLK_IN.n791 CLK_IN.n790 0.00633784
R16654 CLK_IN.n729 CLK_IN.n397 0.00633784
R16655 CLK_IN.n1185 CLK_IN.n45 0.00633784
R16656 CLK_IN.n1263 CLK_IN.n66 0.00633784
R16657 CLK_IN.n967 CLK_IN.n202 0.00590541
R16658 CLK_IN.n1043 CLK_IN.n20 0.00590541
R16659 CLK_IN.n572 CLK_IN.n477 0.00590541
R16660 CLK_IN.n620 CLK_IN.n619 0.00590541
R16661 CLK_IN.n759 CLK_IN.n356 0.00588776
R16662 CLK_IN.n266 CLK_IN.n261 0.00588776
R16663 CLK_IN.n764 CLK_IN.n349 0.00547297
R16664 CLK_IN.n700 CLK_IN.n452 0.00547297
R16665 CLK_IN.n1212 CLK_IN.n54 0.00547297
R16666 CLK_IN.n1291 CLK_IN.n75 0.00547297
R16667 CLK_IN.n794 CLK_IN.n281 0.00525676
R16668 CLK_IN.n731 CLK_IN.n396 0.00525676
R16669 CLK_IN.n1176 CLK_IN.n44 0.00525676
R16670 CLK_IN.n1255 CLK_IN.n65 0.00525676
R16671 CLK_IN.n221 CLK_IN.n215 0.00514865
R16672 CLK_IN.n1067 CLK_IN.n24 0.00514865
R16673 CLK_IN.n558 CLK_IN.n556 0.00514865
R16674 CLK_IN.n629 CLK_IN.n492 0.00514865
R16675 CLK_IN.n1295 CLK_IN.n1294 0.00440238
R16676 CLK_IN.n1000 CLK_IN.n15 0.00439189
R16677 CLK_IN.n599 CLK_IN.n518 0.00439189
R16678 CLK_IN.n822 CLK_IN.n821 0.00439189
R16679 CLK_IN.n359 CLK_IN.n350 0.00439189
R16680 CLK_IN.n1137 CLK_IN.n34 0.00439189
R16681 CLK_IN.n1216 CLK_IN.n55 0.00439189
R16682 CLK_IN.n460 CLK_IN.n459 0.00425921
R16683 CLK_IN.n691 CLK_IN.n461 0.00425921
R16684 CLK_IN.n551 CLK_IN.n548 0.00425921
R16685 CLK_IN.n553 CLK_IN.n529 0.00425921
R16686 CLK_IN.n568 CLK_IN.n526 0.00425921
R16687 CLK_IN.n573 CLK_IN.n570 0.00425921
R16688 CLK_IN.n578 CLK_IN.n524 0.00425921
R16689 CLK_IN.n583 CLK_IN.n522 0.00425921
R16690 CLK_IN.n600 CLK_IN.n597 0.00425921
R16691 CLK_IN.n612 CLK_IN.n609 0.00425921
R16692 CLK_IN.n617 CLK_IN.n514 0.00425921
R16693 CLK_IN.n622 CLK_IN.n512 0.00425921
R16694 CLK_IN.n624 CLK_IN.n511 0.00425921
R16695 CLK_IN.n638 CLK_IN.n636 0.00425921
R16696 CLK_IN.n643 CLK_IN.n507 0.00425921
R16697 CLK_IN.n1300 CLK_IN.n82 0.00425921
R16698 CLK_IN.n90 CLK_IN.n83 0.00425921
R16699 CLK_IN.n324 CLK_IN.n317 0.00425921
R16700 CLK_IN.n783 CLK_IN.n318 0.00425921
R16701 CLK_IN.n424 CLK_IN.n423 0.00425921
R16702 CLK_IN.n719 CLK_IN.n425 0.00425921
R16703 CLK_IN.n1154 CLK_IN.n1153 0.00425921
R16704 CLK_IN.n1159 CLK_IN.n1158 0.00425921
R16705 CLK_IN.n1163 CLK_IN.n1162 0.00425921
R16706 CLK_IN.n1167 CLK_IN.n1166 0.00425921
R16707 CLK_IN.n1188 CLK_IN.n1187 0.00425921
R16708 CLK_IN.n1192 CLK_IN.n1191 0.00425921
R16709 CLK_IN.n1196 CLK_IN.n1195 0.00425921
R16710 CLK_IN.n1200 CLK_IN.n1199 0.00425921
R16711 CLK_IN.n1217 CLK_IN.n1214 0.00425921
R16712 CLK_IN.n1231 CLK_IN.n104 0.00425921
R16713 CLK_IN.n1235 CLK_IN.n1234 0.00425921
R16714 CLK_IN.n1238 CLK_IN.n102 0.00425921
R16715 CLK_IN.n1243 CLK_IN.n100 0.00425921
R16716 CLK_IN.n1266 CLK_IN.n1265 0.00425921
R16717 CLK_IN.n1270 CLK_IN.n1269 0.00425921
R16718 CLK_IN.n1274 CLK_IN.n1273 0.00425921
R16719 CLK_IN.n1277 CLK_IN.n93 0.00425921
R16720 CLK_IN.n442 CLK_IN.n441 0.00424524
R16721 CLK_IN.n536 CLK_IN.n461 0.0042371
R16722 CLK_IN.n540 CLK_IN.n539 0.0042371
R16723 CLK_IN.n544 CLK_IN.n543 0.0042371
R16724 CLK_IN.n548 CLK_IN.n547 0.0042371
R16725 CLK_IN.n559 CLK_IN.n527 0.0042371
R16726 CLK_IN.n564 CLK_IN.n526 0.0042371
R16727 CLK_IN.n584 CLK_IN.n583 0.0042371
R16728 CLK_IN.n588 CLK_IN.n587 0.0042371
R16729 CLK_IN.n592 CLK_IN.n519 0.0042371
R16730 CLK_IN.n597 CLK_IN.n519 0.0042371
R16731 CLK_IN.n601 CLK_IN.n600 0.0042371
R16732 CLK_IN.n605 CLK_IN.n604 0.0042371
R16733 CLK_IN.n609 CLK_IN.n608 0.0042371
R16734 CLK_IN.n628 CLK_IN.n511 0.0042371
R16735 CLK_IN.n631 CLK_IN.n509 0.0042371
R16736 CLK_IN.n645 CLK_IN.n643 0.0042371
R16737 CLK_IN.n650 CLK_IN.n498 0.0042371
R16738 CLK_IN.n505 CLK_IN.n504 0.0042371
R16739 CLK_IN.n501 CLK_IN.n82 0.0042371
R16740 CLK_IN.n289 CLK_IN.n260 0.0042371
R16741 CLK_IN.n797 CLK_IN.n280 0.0042371
R16742 CLK_IN.n311 CLK_IN.n310 0.0042371
R16743 CLK_IN.n353 CLK_IN.n352 0.0042371
R16744 CLK_IN.n751 CLK_IN.n750 0.0042371
R16745 CLK_IN.n406 CLK_IN.n394 0.0042371
R16746 CLK_IN.n732 CLK_IN.n395 0.0042371
R16747 CLK_IN.n706 CLK_IN.n705 0.0042371
R16748 CLK_IN.n456 CLK_IN.n455 0.0042371
R16749 CLK_IN.n1149 CLK_IN.n1148 0.0042371
R16750 CLK_IN.n1153 CLK_IN.n1152 0.0042371
R16751 CLK_IN.n1169 CLK_IN.n1167 0.0042371
R16752 CLK_IN.n1174 CLK_IN.n118 0.0042371
R16753 CLK_IN.n1177 CLK_IN.n116 0.0042371
R16754 CLK_IN.n1187 CLK_IN.n1184 0.0042371
R16755 CLK_IN.n1203 CLK_IN.n1200 0.0042371
R16756 CLK_IN.n1208 CLK_IN.n110 0.0042371
R16757 CLK_IN.n1213 CLK_IN.n108 0.0042371
R16758 CLK_IN.n1214 CLK_IN.n1213 0.0042371
R16759 CLK_IN.n1218 CLK_IN.n1217 0.0042371
R16760 CLK_IN.n1221 CLK_IN.n106 0.0042371
R16761 CLK_IN.n1226 CLK_IN.n104 0.0042371
R16762 CLK_IN.n1248 CLK_IN.n100 0.0042371
R16763 CLK_IN.n1253 CLK_IN.n1250 0.0042371
R16764 CLK_IN.n1256 CLK_IN.n98 0.0042371
R16765 CLK_IN.n1265 CLK_IN.n1262 0.0042371
R16766 CLK_IN.n1282 CLK_IN.n93 0.0042371
R16767 CLK_IN.n1287 CLK_IN.n91 0.0042371
R16768 CLK_IN.n1292 CLK_IN.n1289 0.0042371
R16769 CLK_IN.n1293 CLK_IN.n1292 0.0042371
R16770 CLK_IN.n1141 CLK_IN.n1140 0.00423273
R16771 CLK_IN.n829 CLK_IN.n828 0.00422178
R16772 CLK_IN.n1128 CLK_IN.n133 0.00422178
R16773 CLK_IN.n440 CLK_IN.n422 0.00421905
R16774 CLK_IN.n796 CLK_IN.n278 0.00417568
R16775 CLK_IN.n408 CLK_IN.n407 0.00417568
R16776 CLK_IN.n1172 CLK_IN.n1171 0.00417568
R16777 CLK_IN.n1251 CLK_IN.n64 0.00417568
R16778 CLK_IN.n539 CLK_IN.n535 0.00410442
R16779 CLK_IN.n504 CLK_IN.n499 0.00410442
R16780 CLK_IN.n238 CLK_IN.n233 0.00406757
R16781 CLK_IN.n1097 CLK_IN.n1095 0.00406757
R16782 CLK_IN.n542 CLK_IN.n470 0.00406757
R16783 CLK_IN.n652 CLK_IN.n651 0.00406757
R16784 CLK_IN.n770 CLK_IN.n769 0.00402269
R16785 CLK_IN.n294 CLK_IN.n269 0.00398793
R16786 CLK_IN.n745 CLK_IN.n368 0.00398793
R16787 CLK_IN.n1158 CLK_IN.n122 0.00397174
R16788 CLK_IN.n1196 CLK_IN.n112 0.00397174
R16789 CLK_IN.n1234 CLK_IN.n1232 0.00397174
R16790 CLK_IN.n1278 CLK_IN.n1274 0.00397174
R16791 CLK_IN.n578 CLK_IN.n577 0.00394963
R16792 CLK_IN.n613 CLK_IN.n514 0.00394963
R16793 CLK_IN.n816 CLK_IN.n259 0.00394626
R16794 CLK_IN.n755 CLK_IN.n754 0.00394626
R16795 CLK_IN.n823 CLK_IN.n251 0.00393696
R16796 CLK_IN.n355 CLK_IN.n354 0.00393696
R16797 CLK_IN.n808 CLK_IN.n807 0.00390294
R16798 CLK_IN.n738 CLK_IN.n382 0.00390294
R16799 CLK_IN.n776 CLK_IN.n775 0.00389381
R16800 CLK_IN.n803 CLK_IN.n802 0.00385851
R16801 CLK_IN.n314 CLK_IN.n309 0.00385851
R16802 CLK_IN.n401 CLK_IN.n384 0.00385851
R16803 CLK_IN.n723 CLK_IN.n421 0.00385851
R16804 CLK_IN.n802 CLK_IN.n277 0.00380768
R16805 CLK_IN.n401 CLK_IN.n391 0.00380768
R16806 CLK_IN.n788 CLK_IN.n309 0.00380053
R16807 CLK_IN.n421 CLK_IN.n420 0.00380053
R16808 CLK_IN.n553 CLK_IN.n552 0.00379484
R16809 CLK_IN.n638 CLK_IN.n637 0.00379484
R16810 CLK_IN.n1139 CLK_IN.n132 0.00379484
R16811 CLK_IN.n698 CLK_IN.n457 0.00377273
R16812 CLK_IN.n289 CLK_IN.n267 0.0037725
R16813 CLK_IN.n776 CLK_IN.n337 0.0037725
R16814 CLK_IN.n750 CLK_IN.n365 0.0037725
R16815 CLK_IN.n710 CLK_IN.n709 0.00374762
R16816 CLK_IN.n354 CLK_IN.n351 0.00372958
R16817 CLK_IN.n1168 CLK_IN.n118 0.0037285
R16818 CLK_IN.n1250 CLK_IN.n1249 0.0037285
R16819 CLK_IN.n761 CLK_IN.n353 0.00372177
R16820 CLK_IN.n1183 CLK_IN.n116 0.00370639
R16821 CLK_IN.n1261 CLK_IN.n98 0.00370639
R16822 CLK_IN.n708 CLK_IN.n443 0.00369524
R16823 CLK_IN.n563 CLK_IN.n527 0.00366216
R16824 CLK_IN.n632 CLK_IN.n631 0.00366216
R16825 CLK_IN.n437 CLK_IN.n435 0.00366216
R16826 CLK_IN.n439 CLK_IN.n438 0.00364005
R16827 CLK_IN.n843 CLK_IN.n842 0.00363514
R16828 CLK_IN.n1113 CLK_IN.n30 0.00363514
R16829 CLK_IN.n689 CLK_IN.n463 0.00363514
R16830 CLK_IN.n1302 CLK_IN.n80 0.00363514
R16831 CLK_IN.n1144 CLK_IN.n1142 0.00359048
R16832 CLK_IN.n335 CLK_IN.n318 0.00358532
R16833 CLK_IN.n830 CLK_IN.n829 0.00357902
R16834 CLK_IN.n1128 CLK_IN.n1127 0.00357902
R16835 CLK_IN.n294 CLK_IN.n268 0.00357098
R16836 CLK_IN.n746 CLK_IN.n745 0.00357098
R16837 CLK_IN.n570 CLK_IN.n569 0.00348526
R16838 CLK_IN.n623 CLK_IN.n622 0.00348526
R16839 CLK_IN.n798 CLK_IN.n797 0.003457
R16840 CLK_IN.n406 CLK_IN.n392 0.003457
R16841 CLK_IN.n310 CLK_IN.n308 0.00344926
R16842 CLK_IN.n418 CLK_IN.n395 0.00344926
R16843 CLK_IN.n1163 CLK_IN.n120 0.00344103
R16844 CLK_IN.n1191 CLK_IN.n115 0.00344103
R16845 CLK_IN.n1242 CLK_IN.n102 0.00344103
R16846 CLK_IN.n1269 CLK_IN.n96 0.00344103
R16847 CLK_IN.n322 CLK_IN.n315 0.00343273
R16848 CLK_IN.n724 CLK_IN.n417 0.00343273
R16849 CLK_IN.n804 CLK_IN.n274 0.00341839
R16850 CLK_IN.n737 CLK_IN.n383 0.00341839
R16851 CLK_IN.n390 CLK_IN.n385 0.00341837
R16852 CLK_IN.n812 CLK_IN.n270 0.00341837
R16853 CLK_IN.n1143 CLK_IN.n130 0.00335476
R16854 CLK_IN.n544 CLK_IN.n530 0.00335258
R16855 CLK_IN.n646 CLK_IN.n498 0.00335258
R16856 CLK_IN.n807 CLK_IN.n274 0.0033136
R16857 CLK_IN.n738 CLK_IN.n737 0.0033136
R16858 CLK_IN.n974 CLK_IN.n191 0.00331081
R16859 CLK_IN.n1009 CLK_IN.n16 0.00331081
R16860 CLK_IN.n589 CLK_IN.n481 0.00331081
R16861 CLK_IN.n603 CLK_IN.n485 0.00331081
R16862 CLK_IN.n818 CLK_IN.n257 0.00331081
R16863 CLK_IN.n363 CLK_IN.n361 0.00331081
R16864 CLK_IN.n1147 CLK_IN.n35 0.00331081
R16865 CLK_IN.n1220 CLK_IN.n56 0.00331081
R16866 CLK_IN.n789 CLK_IN.n308 0.00330444
R16867 CLK_IN.n419 CLK_IN.n418 0.00330444
R16868 CLK_IN.n324 CLK_IN.n315 0.0032992
R16869 CLK_IN.n423 CLK_IN.n417 0.0032992
R16870 CLK_IN.n799 CLK_IN.n798 0.00329663
R16871 CLK_IN.n403 CLK_IN.n392 0.00329663
R16872 CLK_IN.n711 CLK_IN.n436 0.00324201
R16873 CLK_IN.n587 CLK_IN.n521 0.00319779
R16874 CLK_IN.n605 CLK_IN.n516 0.00319779
R16875 CLK_IN.n707 CLK_IN.n706 0.00319779
R16876 CLK_IN.n1204 CLK_IN.n110 0.00319779
R16877 CLK_IN.n1281 CLK_IN.n91 0.00319779
R16878 CLK_IN.n816 CLK_IN.n815 0.00317568
R16879 CLK_IN.n754 CLK_IN.n362 0.00317568
R16880 CLK_IN.n1149 CLK_IN.n124 0.00317568
R16881 CLK_IN.n1225 CLK_IN.n106 0.00317568
R16882 CLK_IN.n291 CLK_IN.n268 0.00316007
R16883 CLK_IN.n747 CLK_IN.n746 0.00316007
R16884 CLK_IN.n336 CLK_IN.n335 0.00314581
R16885 CLK_IN.n1145 CLK_IN.n131 0.00310934
R16886 CLK_IN.n801 CLK_IN.n276 0.00309459
R16887 CLK_IN.n402 CLK_IN.n400 0.00309459
R16888 CLK_IN.n119 CLK_IN.n41 0.00309459
R16889 CLK_IN.n1246 CLK_IN.n1245 0.00309459
R16890 CLK_IN.n692 CLK_IN.n460 0.003043
R16891 CLK_IN.n1299 CLK_IN.n83 0.003043
R16892 CLK_IN.n762 CLK_IN.n351 0.00302306
R16893 CLK_IN.n762 CLK_IN.n761 0.00300884
R16894 CLK_IN.n883 CLK_IN.n231 0.0029881
R16895 CLK_IN.n901 CLK_IN.n213 0.0029881
R16896 CLK_IN.n932 CLK_IN.n206 0.0029881
R16897 CLK_IN.n1048 CLK_IN.n1047 0.0029881
R16898 CLK_IN.n337 CLK_IN.n336 0.00298054
R16899 CLK_IN.n291 CLK_IN.n267 0.00298054
R16900 CLK_IN.n747 CLK_IN.n365 0.00298054
R16901 CLK_IN.n1063 CLK_IN.n161 0.0029619
R16902 CLK_IN.n1092 CLK_IN.n1091 0.0029619
R16903 CLK_IN.n789 CLK_IN.n788 0.00293083
R16904 CLK_IN.n420 CLK_IN.n419 0.00293083
R16905 CLK_IN.n799 CLK_IN.n277 0.0029237
R16906 CLK_IN.n403 CLK_IN.n391 0.0029237
R16907 CLK_IN.n593 CLK_IN.n588 0.00291032
R16908 CLK_IN.n604 CLK_IN.n517 0.00291032
R16909 CLK_IN.n769 CLK_IN.n343 0.00291032
R16910 CLK_IN.n705 CLK_IN.n446 0.00291032
R16911 CLK_IN.n1148 CLK_IN.n125 0.00291032
R16912 CLK_IN.n1208 CLK_IN.n1207 0.00291032
R16913 CLK_IN.n1222 CLK_IN.n1221 0.00291032
R16914 CLK_IN.n1288 CLK_IN.n1287 0.00291032
R16915 CLK_IN.n804 CLK_IN.n803 0.00289527
R16916 CLK_IN.n384 CLK_IN.n383 0.00289527
R16917 CLK_IN.n322 CLK_IN.n314 0.00289527
R16918 CLK_IN.n724 CLK_IN.n723 0.00289527
R16919 CLK_IN.n830 CLK_IN.n248 0.00287188
R16920 CLK_IN.n1130 CLK_IN.n1127 0.00284569
R16921 CLK_IN.n775 CLK_IN.n338 0.00283826
R16922 CLK_IN.n1295 CLK_IN.n85 0.00283095
R16923 CLK_IN.n262 CLK_IN.n251 0.00279542
R16924 CLK_IN.n358 CLK_IN.n355 0.00279542
R16925 CLK_IN.n272 CLK_IN.n269 0.00276679
R16926 CLK_IN.n386 CLK_IN.n368 0.00276679
R16927 CLK_IN.n543 CLK_IN.n533 0.00275553
R16928 CLK_IN.n650 CLK_IN.n649 0.00275553
R16929 CLK_IN.n459 CLK_IN.n454 0.00273342
R16930 CLK_IN.n1293 CLK_IN.n90 0.00273342
R16931 CLK_IN.n832 CLK_IN.n248 0.00272619
R16932 CLK_IN.n833 CLK_IN.n832 0.00272619
R16933 CLK_IN.n863 CLK_IN.n862 0.00272619
R16934 CLK_IN.n861 CLK_IN.n839 0.00272619
R16935 CLK_IN.n852 CLK_IN.n851 0.00272619
R16936 CLK_IN.n877 CLK_IN.n876 0.00272619
R16937 CLK_IN.n878 CLK_IN.n877 0.00272619
R16938 CLK_IN.n885 CLK_IN.n884 0.00272619
R16939 CLK_IN.n885 CLK_IN.n227 0.00272619
R16940 CLK_IN.n894 CLK_IN.n225 0.00272619
R16941 CLK_IN.n898 CLK_IN.n225 0.00272619
R16942 CLK_IN.n907 CLK_IN.n906 0.00272619
R16943 CLK_IN.n906 CLK_IN.n900 0.00272619
R16944 CLK_IN.n924 CLK_IN.n923 0.00272619
R16945 CLK_IN.n925 CLK_IN.n924 0.00272619
R16946 CLK_IN.n934 CLK_IN.n931 0.00272619
R16947 CLK_IN.n934 CLK_IN.n933 0.00272619
R16948 CLK_IN.n943 CLK_IN.n942 0.00272619
R16949 CLK_IN.n964 CLK_IN.n963 0.00272619
R16950 CLK_IN.n956 CLK_IN.n955 0.00272619
R16951 CLK_IN.n979 CLK_IN.n196 0.00272619
R16952 CLK_IN.n980 CLK_IN.n979 0.00272619
R16953 CLK_IN.n986 CLK_IN.n985 0.00272619
R16954 CLK_IN.n988 CLK_IN.n986 0.00272619
R16955 CLK_IN.n988 CLK_IN.n987 0.00272619
R16956 CLK_IN.n997 CLK_IN.n996 0.00272619
R16957 CLK_IN.n1006 CLK_IN.n1005 0.00272619
R16958 CLK_IN.n1005 CLK_IN.n182 0.00272619
R16959 CLK_IN.n1015 CLK_IN.n1014 0.00272619
R16960 CLK_IN.n1014 CLK_IN.n179 0.00272619
R16961 CLK_IN.n1021 CLK_IN.n179 0.00272619
R16962 CLK_IN.n1029 CLK_IN.n175 0.00272619
R16963 CLK_IN.n1030 CLK_IN.n1029 0.00272619
R16964 CLK_IN.n1039 CLK_IN.n1038 0.00272619
R16965 CLK_IN.n1040 CLK_IN.n1039 0.00272619
R16966 CLK_IN.n1053 CLK_IN.n169 0.00272619
R16967 CLK_IN.n1062 CLK_IN.n1061 0.00272619
R16968 CLK_IN.n1070 CLK_IN.n1069 0.00272619
R16969 CLK_IN.n1072 CLK_IN.n1071 0.00272619
R16970 CLK_IN.n1080 CLK_IN.n153 0.00272619
R16971 CLK_IN.n1090 CLK_IN.n1089 0.00272619
R16972 CLK_IN.n1092 CLK_IN.n1090 0.00272619
R16973 CLK_IN.n1100 CLK_IN.n147 0.00272619
R16974 CLK_IN.n1101 CLK_IN.n1100 0.00272619
R16975 CLK_IN.n1102 CLK_IN.n1101 0.00272619
R16976 CLK_IN.n1110 CLK_IN.n1108 0.00272619
R16977 CLK_IN.n1110 CLK_IN.n1109 0.00272619
R16978 CLK_IN.n1119 CLK_IN.n1117 0.00272619
R16979 CLK_IN.n1119 CLK_IN.n1118 0.00272619
R16980 CLK_IN.n1133 CLK_IN.n1132 0.00272619
R16981 CLK_IN.n1131 CLK_IN.n1130 0.00272619
R16982 CLK_IN.n833 CLK_IN.n246 0.0027
R16983 CLK_IN.n862 CLK_IN.n861 0.0027
R16984 CLK_IN.n852 CLK_IN.n841 0.0027
R16985 CLK_IN.n876 CLK_IN.n234 0.0027
R16986 CLK_IN.n884 CLK_IN.n883 0.0027
R16987 CLK_IN.n902 CLK_IN.n900 0.0027
R16988 CLK_IN.n964 CLK_IN.n943 0.0027
R16989 CLK_IN.n957 CLK_IN.n956 0.0027
R16990 CLK_IN.n949 CLK_IN.n196 0.0027
R16991 CLK_IN.n997 CLK_IN.n995 0.0027
R16992 CLK_IN.n1006 CLK_IN.n1004 0.0027
R16993 CLK_IN.n1040 CLK_IN.n171 0.0027
R16994 CLK_IN.n1049 CLK_IN.n169 0.0027
R16995 CLK_IN.n1061 CLK_IN.n165 0.0027
R16996 CLK_IN.n1072 CLK_IN.n1070 0.0027
R16997 CLK_IN.n1080 CLK_IN.n1079 0.0027
R16998 CLK_IN.n1089 CLK_IN.n151 0.0027
R16999 CLK_IN.n1118 CLK_IN.n137 0.0027
R17000 CLK_IN.n1132 CLK_IN.n1131 0.0027
R17001 CLK_IN.n902 CLK_IN.n901 0.00264762
R17002 CLK_IN.n1069 CLK_IN.n161 0.00264762
R17003 CLK_IN.n1162 CLK_IN.n121 0.00264496
R17004 CLK_IN.n1239 CLK_IN.n1238 0.00264496
R17005 CLK_IN.n784 CLK_IN.n317 0.00262285
R17006 CLK_IN.n720 CLK_IN.n424 0.00262285
R17007 CLK_IN.n1192 CLK_IN.n113 0.00262285
R17008 CLK_IN.n1270 CLK_IN.n95 0.00262285
R17009 CLK_IN.n933 CLK_IN.n932 0.00262143
R17010 CLK_IN.n1049 CLK_IN.n1048 0.00262143
R17011 CLK_IN.n574 CLK_IN.n573 0.00260074
R17012 CLK_IN.n616 CLK_IN.n512 0.00260074
R17013 CLK_IN.n881 CLK_IN.n880 0.00257862
R17014 CLK_IN.n1093 CLK_IN.n148 0.00257862
R17015 CLK_IN.n1047 CLK_IN.n171 0.00256905
R17016 CLK_IN.n937 CLK_IN.n936 0.00255405
R17017 CLK_IN.n167 CLK_IN.n21 0.00255405
R17018 CLK_IN.n567 CLK_IN.n476 0.00255405
R17019 CLK_IN.n625 CLK_IN.n490 0.00255405
R17020 CLK_IN.n942 CLK_IN.n206 0.00254286
R17021 CLK_IN.n1063 CLK_IN.n1062 0.00254286
R17022 CLK_IN.n940 CLK_IN.n939 0.0025344
R17023 CLK_IN.n923 CLK_IN.n213 0.00251667
R17024 CLK_IN.n1046 CLK_IN.n1045 0.00251228
R17025 CLK_IN.n827 CLK_IN.n826 0.0024936
R17026 CLK_IN.n878 CLK_IN.n231 0.00246429
R17027 CLK_IN.n1091 CLK_IN.n147 0.00246429
R17028 CLK_IN.n560 CLK_IN.n559 0.00244595
R17029 CLK_IN.n635 CLK_IN.n509 0.00244595
R17030 CLK_IN.n899 CLK_IN.n898 0.0024381
R17031 CLK_IN.n1079 CLK_IN.n1078 0.0024381
R17032 CLK_IN.n920 CLK_IN.n214 0.00242383
R17033 CLK_IN.n1065 CLK_IN.n162 0.00242383
R17034 CLK_IN.n1142 CLK_IN.n1141 0.00238571
R17035 CLK_IN.n710 CLK_IN.n442 0.00238571
R17036 CLK_IN.n857 CLK_IN.n856 0.00238571
R17037 CLK_IN.n850 CLK_IN.n846 0.00238571
R17038 CLK_IN.n893 CLK_IN.n892 0.00238571
R17039 CLK_IN.n908 CLK_IN.n899 0.00238571
R17040 CLK_IN.n930 CLK_IN.n211 0.00238571
R17041 CLK_IN.n962 CLK_IN.n944 0.00238571
R17042 CLK_IN.n950 CLK_IN.n948 0.00238571
R17043 CLK_IN.n994 CLK_IN.n189 0.00238571
R17044 CLK_IN.n1003 CLK_IN.n185 0.00238571
R17045 CLK_IN.n1012 CLK_IN.n182 0.00238571
R17046 CLK_IN.n1023 CLK_IN.n1022 0.00238571
R17047 CLK_IN.n1031 CLK_IN.n173 0.00238571
R17048 CLK_IN.n1055 CLK_IN.n1054 0.00238571
R17049 CLK_IN.n1078 CLK_IN.n157 0.00238571
R17050 CLK_IN.n1085 CLK_IN.n1084 0.00238571
R17051 CLK_IN.n1107 CLK_IN.n145 0.00238571
R17052 CLK_IN.n1116 CLK_IN.n140 0.00238571
R17053 CLK_IN.n864 CLK_IN.n245 0.00237961
R17054 CLK_IN.n860 CLK_IN.n859 0.00237961
R17055 CLK_IN.n853 CLK_IN.n845 0.00237961
R17056 CLK_IN.n875 CLK_IN.n232 0.00237961
R17057 CLK_IN.n879 CLK_IN.n232 0.00237961
R17058 CLK_IN.n886 CLK_IN.n230 0.00237961
R17059 CLK_IN.n886 CLK_IN.n228 0.00237961
R17060 CLK_IN.n896 CLK_IN.n895 0.00237961
R17061 CLK_IN.n897 CLK_IN.n896 0.00237961
R17062 CLK_IN.n905 CLK_IN.n224 0.00237961
R17063 CLK_IN.n905 CLK_IN.n904 0.00237961
R17064 CLK_IN.n922 CLK_IN.n212 0.00237961
R17065 CLK_IN.n926 CLK_IN.n212 0.00237961
R17066 CLK_IN.n935 CLK_IN.n209 0.00237961
R17067 CLK_IN.n935 CLK_IN.n210 0.00237961
R17068 CLK_IN.n941 CLK_IN.n204 0.00237961
R17069 CLK_IN.n965 CLK_IN.n205 0.00237961
R17070 CLK_IN.n954 CLK_IN.n947 0.00237961
R17071 CLK_IN.n978 CLK_IN.n977 0.00237961
R17072 CLK_IN.n978 CLK_IN.n195 0.00237961
R17073 CLK_IN.n984 CLK_IN.n192 0.00237961
R17074 CLK_IN.n989 CLK_IN.n192 0.00237961
R17075 CLK_IN.n989 CLK_IN.n193 0.00237961
R17076 CLK_IN.n998 CLK_IN.n188 0.00237961
R17077 CLK_IN.n1007 CLK_IN.n183 0.00237961
R17078 CLK_IN.n1010 CLK_IN.n183 0.00237961
R17079 CLK_IN.n1016 CLK_IN.n180 0.00237961
R17080 CLK_IN.n1019 CLK_IN.n180 0.00237961
R17081 CLK_IN.n1020 CLK_IN.n1019 0.00237961
R17082 CLK_IN.n1028 CLK_IN.n176 0.00237961
R17083 CLK_IN.n1028 CLK_IN.n174 0.00237961
R17084 CLK_IN.n1037 CLK_IN.n172 0.00237961
R17085 CLK_IN.n1041 CLK_IN.n172 0.00237961
R17086 CLK_IN.n1052 CLK_IN.n1051 0.00237961
R17087 CLK_IN.n1060 CLK_IN.n164 0.00237961
R17088 CLK_IN.n1068 CLK_IN.n159 0.00237961
R17089 CLK_IN.n1073 CLK_IN.n160 0.00237961
R17090 CLK_IN.n1082 CLK_IN.n1081 0.00237961
R17091 CLK_IN.n1088 CLK_IN.n150 0.00237961
R17092 CLK_IN.n1093 CLK_IN.n150 0.00237961
R17093 CLK_IN.n1099 CLK_IN.n1098 0.00237961
R17094 CLK_IN.n1099 CLK_IN.n146 0.00237961
R17095 CLK_IN.n1103 CLK_IN.n146 0.00237961
R17096 CLK_IN.n1111 CLK_IN.n143 0.00237961
R17097 CLK_IN.n1111 CLK_IN.n144 0.00237961
R17098 CLK_IN.n1120 CLK_IN.n139 0.00237961
R17099 CLK_IN.n1120 CLK_IN.n138 0.00237961
R17100 CLK_IN.n1134 CLK_IN.n134 0.00237961
R17101 CLK_IN.n825 CLK_IN.n247 0.00237961
R17102 CLK_IN.n264 CLK_IN.n263 0.00237961
R17103 CLK_IN.n312 CLK_IN.n280 0.00237961
R17104 CLK_IN.n312 CLK_IN.n311 0.00237961
R17105 CLK_IN.n772 CLK_IN.n771 0.00237961
R17106 CLK_IN.n757 CLK_IN.n756 0.00237961
R17107 CLK_IN.n733 CLK_IN.n394 0.00237961
R17108 CLK_IN.n733 CLK_IN.n732 0.00237961
R17109 CLK_IN.n1178 CLK_IN.n1174 0.00237961
R17110 CLK_IN.n1178 CLK_IN.n1177 0.00237961
R17111 CLK_IN.n1257 CLK_IN.n1253 0.00237961
R17112 CLK_IN.n1257 CLK_IN.n1256 0.00237961
R17113 CLK_IN.n957 CLK_IN.n944 0.00235952
R17114 CLK_IN.n985 CLK_IN.n194 0.00235952
R17115 CLK_IN.n835 CLK_IN.n834 0.00235749
R17116 CLK_IN.n860 CLK_IN.n245 0.00235749
R17117 CLK_IN.n854 CLK_IN.n853 0.00235749
R17118 CLK_IN.n875 CLK_IN.n235 0.00235749
R17119 CLK_IN.n882 CLK_IN.n230 0.00235749
R17120 CLK_IN.n904 CLK_IN.n903 0.00235749
R17121 CLK_IN.n965 CLK_IN.n204 0.00235749
R17122 CLK_IN.n958 CLK_IN.n947 0.00235749
R17123 CLK_IN.n977 CLK_IN.n197 0.00235749
R17124 CLK_IN.n998 CLK_IN.n187 0.00235749
R17125 CLK_IN.n1007 CLK_IN.n184 0.00235749
R17126 CLK_IN.n1042 CLK_IN.n1041 0.00235749
R17127 CLK_IN.n1051 CLK_IN.n1050 0.00235749
R17128 CLK_IN.n1060 CLK_IN.n166 0.00235749
R17129 CLK_IN.n1073 CLK_IN.n159 0.00235749
R17130 CLK_IN.n1081 CLK_IN.n154 0.00235749
R17131 CLK_IN.n1088 CLK_IN.n1087 0.00235749
R17132 CLK_IN.n1123 CLK_IN.n138 0.00235749
R17133 CLK_IN.n810 CLK_IN.n809 0.00235749
R17134 CLK_IN.n388 CLK_IN.n387 0.00235749
R17135 CLK_IN.n1031 CLK_IN.n1030 0.00233333
R17136 CLK_IN.n903 CLK_IN.n214 0.00231327
R17137 CLK_IN.n1068 CLK_IN.n162 0.00231327
R17138 CLK_IN.n837 CLK_IN.n246 0.00230714
R17139 CLK_IN.n1125 CLK_IN.n137 0.00230714
R17140 CLK_IN.n1133 CLK_IN.n1126 0.00230714
R17141 CLK_IN.n210 CLK_IN.n207 0.00229115
R17142 CLK_IN.n1050 CLK_IN.n170 0.00229115
R17143 CLK_IN.n560 CLK_IN.n529 0.00229115
R17144 CLK_IN.n636 CLK_IN.n635 0.00229115
R17145 CLK_IN.n863 CLK_IN.n838 0.00228095
R17146 CLK_IN.n851 CLK_IN.n850 0.00228095
R17147 CLK_IN.n1108 CLK_IN.n1107 0.00225476
R17148 CLK_IN.n1046 CLK_IN.n1042 0.00224693
R17149 CLK_IN.n288 CLK_IN.n258 0.00222973
R17150 CLK_IN.n752 CLK_IN.n364 0.00222973
R17151 CLK_IN.n1151 CLK_IN.n36 0.00222973
R17152 CLK_IN.n1228 CLK_IN.n1227 0.00222973
R17153 CLK_IN.n941 CLK_IN.n940 0.00222482
R17154 CLK_IN.n1064 CLK_IN.n164 0.00222482
R17155 CLK_IN.n922 CLK_IN.n921 0.0022027
R17156 CLK_IN.n981 CLK_IN.n980 0.00220238
R17157 CLK_IN.n1015 CLK_IN.n1013 0.00220238
R17158 CLK_IN.n995 CLK_IN.n994 0.00217619
R17159 CLK_IN.n996 CLK_IN.n185 0.00217619
R17160 CLK_IN.n880 CLK_IN.n879 0.00215848
R17161 CLK_IN.n1098 CLK_IN.n148 0.00215848
R17162 CLK_IN.n897 CLK_IN.n223 0.00213636
R17163 CLK_IN.n1077 CLK_IN.n154 0.00213636
R17164 CLK_IN.n574 CLK_IN.n524 0.00213636
R17165 CLK_IN.n617 CLK_IN.n616 0.00213636
R17166 CLK_IN.n784 CLK_IN.n783 0.00211425
R17167 CLK_IN.n720 CLK_IN.n719 0.00211425
R17168 CLK_IN.n1195 CLK_IN.n113 0.00211425
R17169 CLK_IN.n1273 CLK_IN.n95 0.00211425
R17170 CLK_IN.n1144 CLK_IN.n1143 0.00209762
R17171 CLK_IN.n856 CLK_IN.n841 0.00209762
R17172 CLK_IN.n1011 CLK_IN.n1010 0.00209214
R17173 CLK_IN.n811 CLK_IN.n272 0.00209214
R17174 CLK_IN.n389 CLK_IN.n386 0.00209214
R17175 CLK_IN.n1159 CLK_IN.n121 0.00209214
R17176 CLK_IN.n1239 CLK_IN.n1235 0.00209214
R17177 CLK_IN.n1109 CLK_IN.n140 0.00207143
R17178 CLK_IN.n959 CLK_IN.n958 0.00207002
R17179 CLK_IN.n984 CLK_IN.n983 0.00207002
R17180 CLK_IN.n1032 CLK_IN.n174 0.00204791
R17181 CLK_IN.n836 CLK_IN.n835 0.0020258
R17182 CLK_IN.n1124 CLK_IN.n1123 0.0020258
R17183 CLK_IN.n1134 CLK_IN.n136 0.0020258
R17184 CLK_IN.n955 CLK_IN.n948 0.00201905
R17185 CLK_IN.n806 CLK_IN.n275 0.00201351
R17186 CLK_IN.n740 CLK_IN.n739 0.00201351
R17187 CLK_IN.n1164 CLK_IN.n40 0.00201351
R17188 CLK_IN.n101 CLK_IN.n61 0.00201351
R17189 CLK_IN.n864 CLK_IN.n244 0.00200369
R17190 CLK_IN.n849 CLK_IN.n845 0.00200369
R17191 CLK_IN.n540 CLK_IN.n533 0.00200369
R17192 CLK_IN.n649 CLK_IN.n505 0.00200369
R17193 CLK_IN.n828 CLK_IN.n827 0.00200107
R17194 CLK_IN.n826 CLK_IN.n250 0.00200107
R17195 CLK_IN.n1140 CLK_IN.n133 0.00200107
R17196 CLK_IN.n1023 CLK_IN.n175 0.00199286
R17197 CLK_IN.n1106 CLK_IN.n143 0.00198157
R17198 CLK_IN.n982 CLK_IN.n195 0.00193735
R17199 CLK_IN.n1016 CLK_IN.n181 0.00193735
R17200 CLK_IN.n993 CLK_IN.n187 0.00191523
R17201 CLK_IN.n188 CLK_IN.n186 0.00191523
R17202 CLK_IN.n831 CLK_IN.n247 0.00191523
R17203 CLK_IN.n825 CLK_IN.n824 0.00191523
R17204 CLK_IN.n1139 CLK_IN.n135 0.00191523
R17205 CLK_IN.n1293 CLK_IN.n86 0.00191523
R17206 CLK_IN.n894 CLK_IN.n893 0.00191429
R17207 CLK_IN.n1084 CLK_IN.n153 0.00191429
R17208 CLK_IN.n910 CLK_IN.n909 0.00187101
R17209 CLK_IN.n809 CLK_IN.n808 0.00185493
R17210 CLK_IN.n387 CLK_IN.n382 0.00185493
R17211 CLK_IN.n855 CLK_IN.n854 0.00184889
R17212 CLK_IN.n1076 CLK_IN.n158 0.00184889
R17213 CLK_IN.n593 CLK_IN.n592 0.00184889
R17214 CLK_IN.n601 CLK_IN.n517 0.00184889
R17215 CLK_IN.n265 CLK_IN.n262 0.00184889
R17216 CLK_IN.n352 CLK_IN.n343 0.00184889
R17217 CLK_IN.n758 CLK_IN.n358 0.00184889
R17218 CLK_IN.n455 CLK_IN.n446 0.00184889
R17219 CLK_IN.n1145 CLK_IN.n125 0.00184889
R17220 CLK_IN.n1207 CLK_IN.n108 0.00184889
R17221 CLK_IN.n1222 CLK_IN.n1218 0.00184889
R17222 CLK_IN.n1289 CLK_IN.n1288 0.00184889
R17223 CLK_IN.n1055 CLK_IN.n165 0.00183571
R17224 CLK_IN.n144 CLK_IN.n141 0.00182678
R17225 CLK_IN.n925 CLK_IN.n211 0.00180952
R17226 CLK_IN.n918 CLK_IN.n216 0.0017973
R17227 CLK_IN.n1059 CLK_IN.n163 0.0017973
R17228 CLK_IN.n565 CLK_IN.n475 0.0017973
R17229 CLK_IN.n627 CLK_IN.n491 0.0017973
R17230 CLK_IN.n263 CLK_IN.n259 0.0017897
R17231 CLK_IN.n756 CLK_IN.n755 0.0017897
R17232 CLK_IN.n961 CLK_IN.n960 0.00178256
R17233 CLK_IN.n954 CLK_IN.n953 0.00178256
R17234 CLK_IN.n1036 CLK_IN.n1035 0.00178256
R17235 CLK_IN.n1024 CLK_IN.n176 0.00176044
R17236 CLK_IN.n709 CLK_IN.n708 0.00175714
R17237 CLK_IN.n931 CLK_IN.n930 0.00173095
R17238 CLK_IN.n1054 CLK_IN.n1053 0.00173095
R17239 CLK_IN.n848 CLK_IN.n847 0.00171622
R17240 CLK_IN.n771 CLK_IN.n770 0.00171347
R17241 CLK_IN.n895 CLK_IN.n226 0.0016941
R17242 CLK_IN.n1083 CLK_IN.n1082 0.0016941
R17243 CLK_IN.n1105 CLK_IN.n1104 0.0016941
R17244 CLK_IN.n692 CLK_IN.n691 0.0016941
R17245 CLK_IN.n1300 CLK_IN.n1299 0.0016941
R17246 CLK_IN.n1085 CLK_IN.n151 0.00165238
R17247 CLK_IN.n992 CLK_IN.n190 0.00162776
R17248 CLK_IN.n1002 CLK_IN.n1001 0.00162776
R17249 CLK_IN.n1056 CLK_IN.n166 0.00162776
R17250 CLK_IN.n1136 CLK_IN.n131 0.00162776
R17251 CLK_IN.n892 CLK_IN.n227 0.00162619
R17252 CLK_IN.n927 CLK_IN.n926 0.00160565
R17253 CLK_IN.n815 CLK_IN.n260 0.00158354
R17254 CLK_IN.n751 CLK_IN.n362 0.00158354
R17255 CLK_IN.n1152 CLK_IN.n124 0.00158354
R17256 CLK_IN.n1226 CLK_IN.n1225 0.00158354
R17257 CLK_IN.n858 CLK_IN.n840 0.00156143
R17258 CLK_IN.n1115 CLK_IN.n1114 0.00156143
R17259 CLK_IN.n584 CLK_IN.n521 0.00156143
R17260 CLK_IN.n608 CLK_IN.n516 0.00156143
R17261 CLK_IN.n773 CLK_IN.n338 0.00156143
R17262 CLK_IN.n707 CLK_IN.n436 0.00156143
R17263 CLK_IN.n1204 CLK_IN.n1203 0.00156143
R17264 CLK_IN.n1282 CLK_IN.n1281 0.00156143
R17265 CLK_IN.n950 CLK_IN.n949 0.00154762
R17266 CLK_IN.n1022 CLK_IN.n1021 0.00154762
R17267 CLK_IN.n929 CLK_IN.n209 0.00153931
R17268 CLK_IN.n1052 CLK_IN.n168 0.00153931
R17269 CLK_IN.n952 CLK_IN.n951 0.00149509
R17270 CLK_IN.n712 CLK_IN.n711 0.00149509
R17271 CLK_IN.n1025 CLK_IN.n178 0.00147297
R17272 CLK_IN.n1087 CLK_IN.n1086 0.00147297
R17273 CLK_IN.n857 CLK_IN.n839 0.00146905
R17274 CLK_IN.n1117 CLK_IN.n1116 0.00146905
R17275 CLK_IN.n891 CLK_IN.n228 0.00145086
R17276 CLK_IN.n891 CLK_IN.n890 0.00140663
R17277 CLK_IN.n1086 CLK_IN.n152 0.00140663
R17278 CLK_IN.n547 CLK_IN.n530 0.00140663
R17279 CLK_IN.n646 CLK_IN.n645 0.00140663
R17280 CLK_IN.n1004 CLK_IN.n1003 0.00139048
R17281 CLK_IN.n951 CLK_IN.n197 0.00138452
R17282 CLK_IN.n1020 CLK_IN.n178 0.00138452
R17283 CLK_IN.n838 CLK_IN.n837 0.00136429
R17284 CLK_IN.n981 CLK_IN.n194 0.00136429
R17285 CLK_IN.n987 CLK_IN.n189 0.00136429
R17286 CLK_IN.n929 CLK_IN.n928 0.00134029
R17287 CLK_IN.n1057 CLK_IN.n168 0.00134029
R17288 CLK_IN.n1013 CLK_IN.n1012 0.00133809
R17289 CLK_IN.n1126 CLK_IN.n1125 0.00133809
R17290 CLK_IN.n859 CLK_IN.n858 0.00131818
R17291 CLK_IN.n1115 CLK_IN.n139 0.00131818
R17292 CLK_IN.n773 CLK_IN.n772 0.00131818
R17293 CLK_IN.n1166 CLK_IN.n120 0.00129607
R17294 CLK_IN.n1188 CLK_IN.n115 0.00129607
R17295 CLK_IN.n1243 CLK_IN.n1242 0.00129607
R17296 CLK_IN.n1266 CLK_IN.n96 0.00129607
R17297 CLK_IN.n846 CLK_IN.n234 0.00128571
R17298 CLK_IN.n1102 CLK_IN.n145 0.00128571
R17299 CLK_IN.n928 CLK_IN.n927 0.00125184
R17300 CLK_IN.n1002 CLK_IN.n184 0.00125184
R17301 CLK_IN.n1057 CLK_IN.n1056 0.00125184
R17302 CLK_IN.n569 CLK_IN.n568 0.00125184
R17303 CLK_IN.n624 CLK_IN.n623 0.00125184
R17304 CLK_IN.n836 CLK_IN.n244 0.00122973
R17305 CLK_IN.n983 CLK_IN.n982 0.00122973
R17306 CLK_IN.n193 CLK_IN.n190 0.00122973
R17307 CLK_IN.n1011 CLK_IN.n181 0.00120762
R17308 CLK_IN.n1124 CLK_IN.n136 0.00120762
R17309 CLK_IN.n963 CLK_IN.n962 0.00120714
R17310 CLK_IN.n1038 CLK_IN.n173 0.00120714
R17311 CLK_IN.n890 CLK_IN.n226 0.0011855
R17312 CLK_IN.n1083 CLK_IN.n152 0.0011855
R17313 CLK_IN.n847 CLK_IN.n235 0.00116339
R17314 CLK_IN.n1104 CLK_IN.n1103 0.00116339
R17315 CLK_IN.n293 CLK_IN.n292 0.00114865
R17316 CLK_IN.n748 CLK_IN.n366 0.00114865
R17317 CLK_IN.n1156 CLK_IN.n1155 0.00114865
R17318 CLK_IN.n1230 CLK_IN.n59 0.00114865
R17319 CLK_IN.n1071 CLK_IN.n157 0.00112857
R17320 CLK_IN.n1025 CLK_IN.n1024 0.00111916
R17321 CLK_IN.n908 CLK_IN.n907 0.00110238
R17322 CLK_IN.n961 CLK_IN.n205 0.00109705
R17323 CLK_IN.n953 CLK_IN.n952 0.00109705
R17324 CLK_IN.n1037 CLK_IN.n1036 0.00109705
R17325 CLK_IN.n564 CLK_IN.n563 0.00109705
R17326 CLK_IN.n632 CLK_IN.n628 0.00109705
R17327 CLK_IN.n712 CLK_IN.n435 0.00109705
R17328 CLK_IN.n1184 CLK_IN.n1183 0.00105283
R17329 CLK_IN.n1262 CLK_IN.n1261 0.00105283
R17330 CLK_IN.n1296 CLK_IN.n86 0.00105283
R17331 CLK_IN.n991 CLK_IN.n14 0.00104054
R17332 CLK_IN.n590 CLK_IN.n482 0.00104054
R17333 CLK_IN.n855 CLK_IN.n840 0.00103071
R17334 CLK_IN.n160 CLK_IN.n158 0.00103071
R17335 CLK_IN.n1114 CLK_IN.n141 0.00103071
R17336 CLK_IN.n831 CLK_IN.n249 0.00103071
R17337 CLK_IN.n265 CLK_IN.n264 0.00103071
R17338 CLK_IN.n758 CLK_IN.n757 0.00103071
R17339 CLK_IN.n1129 CLK_IN.n135 0.00103071
R17340 CLK_IN.n1169 CLK_IN.n1168 0.00103071
R17341 CLK_IN.n1249 CLK_IN.n1248 0.00103071
R17342 CLK_IN.n909 CLK_IN.n224 0.0010086
R17343 CLK_IN.n993 CLK_IN.n992 0.000964373
R17344 CLK_IN.n1001 CLK_IN.n186 0.000964373
R17345 CLK_IN.n824 CLK_IN.n823 0.000964373
R17346 CLK_IN.n457 CLK_IN.n456 0.000964373
R17347 CLK_IN.n1136 CLK_IN.n132 0.000964373
R17348 CLK_IN.n552 CLK_IN.n551 0.00094226
R17349 CLK_IN.n637 CLK_IN.n507 0.00094226
R17350 CLK_IN.n297 CLK_IN.n296 0.000932432
R17351 CLK_IN.n743 CLK_IN.n369 0.000932432
R17352 CLK_IN.n1160 CLK_IN.n39 0.000932432
R17353 CLK_IN.n1236 CLK_IN.n60 0.000932432
R17354 CLK_IN.n834 CLK_IN.n247 0.000898034
R17355 CLK_IN.n1106 CLK_IN.n1105 0.000898034
R17356 CLK_IN.n849 CLK_IN.n848 0.000875921
R17357 CLK_IN.n1139 CLK_IN.n134 0.000853808
R17358 CLK_IN.n438 CLK_IN.n425 0.000831695
R17359 CLK_IN.n441 CLK_IN.n440 0.000814286
R17360 CLK_IN.n960 CLK_IN.n959 0.000809582
R17361 CLK_IN.n1035 CLK_IN.n1032 0.000809582
R17362 CLK_IN.n577 CLK_IN.n522 0.000787469
R17363 CLK_IN.n613 CLK_IN.n612 0.000787469
R17364 CLK_IN.n811 CLK_IN.n810 0.000787469
R17365 CLK_IN.n389 CLK_IN.n388 0.000787469
R17366 CLK_IN.n439 CLK_IN.n437 0.000765356
R17367 CLK_IN.n1154 CLK_IN.n122 0.000765356
R17368 CLK_IN.n1199 CLK_IN.n112 0.000765356
R17369 CLK_IN.n1232 CLK_IN.n1231 0.000765356
R17370 CLK_IN.n1278 CLK_IN.n1277 0.000765356
R17371 CLK_IN.n1077 CLK_IN.n1076 0.000743243
R17372 CLK_IN.n910 CLK_IN.n223 0.00072113
R17373 CLK_IN.n873 CLK_IN.n236 0.000716216
R17374 CLK_IN.n142 CLK_IN.n29 0.000716216
R17375 CLK_IN.n538 CLK_IN.n534 0.000716216
R17376 CLK_IN.n503 CLK_IN.n500 0.000716216
R17377 CLK_IN.n921 CLK_IN.n920 0.000676904
R17378 CLK_IN.n1065 CLK_IN.n1064 0.000654791
R17379 CLK_IN.n536 CLK_IN.n535 0.000654791
R17380 CLK_IN.n501 CLK_IN.n499 0.000654791
R17381 CLK_IN.n1045 CLK_IN.n170 0.000588452
R17382 CLK_IN.n939 CLK_IN.n207 0.000566339
R17383 CLK_IN.n882 CLK_IN.n881 0.000522113
R17384 CLK_IN.n698 CLK_IN.n454 0.000522113
R17385 X0.n3 X0.n0 15.1893
R17386 X0.n2 X0.n1 15.0005
R17387 X0 X0.n3 9.55138
R17388 X0.n897 X0.n280 2.2505
R17389 X0.n895 X0.n282 2.2505
R17390 X0.n891 X0.n285 2.2505
R17391 X0.n889 X0.n287 2.2505
R17392 X0.n885 X0.n884 2.2505
R17393 X0.n1374 X0.n7 2.2505
R17394 X0.n1372 X0.n9 2.2505
R17395 X0.n1368 X0.n12 2.2505
R17396 X0.n1367 X0.n13 2.2505
R17397 X0.n462 X0.n15 2.2505
R17398 X0.n1361 X0.n18 2.2505
R17399 X0.n483 X0.n20 2.2505
R17400 X0.n1355 X0.n23 2.2505
R17401 X0.n504 X0.n25 2.2505
R17402 X0.n1349 X0.n28 2.2505
R17403 X0.n1284 X0.n73 2.2505
R17404 X0.n89 X0.n82 2.2505
R17405 X0.n1266 X0.n84 2.2505
R17406 X0.n1258 X0.n1257 2.2505
R17407 X0.n1252 X0.n1251 2.2505
R17408 X0.n116 X0.n112 2.2505
R17409 X0.n1208 X0.n115 2.2505
R17410 X0.n1219 X0.n1218 2.2505
R17411 X0.n1196 X0.n1195 2.2505
R17412 X0.n1191 X0.n1190 2.2505
R17413 X0.n1156 X0.n137 2.2505
R17414 X0.n1161 X0.n1160 2.2505
R17415 X0.n1153 X0.n1152 2.2505
R17416 X0.n1134 X0.n1133 2.2505
R17417 X0.n1129 X0.n1128 2.2505
R17418 X0.n1279 X0.n73 2.2505
R17419 X0.n1278 X0.n82 2.2505
R17420 X0.n84 X0.n83 2.2505
R17421 X0.n1257 X0.n1256 2.2505
R17422 X0.n1253 X0.n1252 2.2505
R17423 X0.n1222 X0.n116 2.2505
R17424 X0.n1221 X0.n115 2.2505
R17425 X0.n1220 X0.n1219 2.2505
R17426 X0.n1195 X0.n1194 2.2505
R17427 X0.n1192 X0.n1191 2.2505
R17428 X0.n1157 X0.n1156 2.2505
R17429 X0.n1160 X0.n1159 2.2505
R17430 X0.n1154 X0.n1153 2.2505
R17431 X0.n1133 X0.n1132 2.2505
R17432 X0.n1130 X0.n1129 2.2505
R17433 X0.n1118 X0.n1117 2.2505
R17434 X0.n1116 X0.n171 2.2505
R17435 X0.n1115 X0.n1114 2.2505
R17436 X0.n173 X0.n172 2.2505
R17437 X0.n1087 X0.n1086 2.2505
R17438 X0.n1085 X0.n185 2.2505
R17439 X0.n1084 X0.n1083 2.2505
R17440 X0.n187 X0.n186 2.2505
R17441 X0.n1061 X0.n1060 2.2505
R17442 X0.n1059 X0.n198 2.2505
R17443 X0.n1058 X0.n1057 2.2505
R17444 X0.n200 X0.n199 2.2505
R17445 X0.n1022 X0.n1021 2.2505
R17446 X0.n1029 X0.n1020 2.2505
R17447 X0.n1030 X0.n1019 2.2505
R17448 X0.n1018 X0.n216 2.2505
R17449 X0.n1017 X0.n1016 2.2505
R17450 X0.n218 X0.n217 2.2505
R17451 X0.n1000 X0.n999 2.2505
R17452 X0.n998 X0.n233 2.2505
R17453 X0.n997 X0.n996 2.2505
R17454 X0.n235 X0.n234 2.2505
R17455 X0.n956 X0.n955 2.2505
R17456 X0.n963 X0.n954 2.2505
R17457 X0.n964 X0.n953 2.2505
R17458 X0.n952 X0.n252 2.2505
R17459 X0.n951 X0.n950 2.2505
R17460 X0.n254 X0.n253 2.2505
R17461 X0.n929 X0.n928 2.2505
R17462 X0.n927 X0.n265 2.2505
R17463 X0.n926 X0.n925 2.2505
R17464 X0.n267 X0.n266 2.2505
R17465 X0.n902 X0.n901 2.2505
R17466 X0.n903 X0.n900 2.2505
R17467 X0.n904 X0.n903 2.2505
R17468 X0.n902 X0.n271 2.2505
R17469 X0.n916 X0.n267 2.2505
R17470 X0.n925 X0.n924 2.2505
R17471 X0.n269 X0.n265 2.2505
R17472 X0.n930 X0.n929 2.2505
R17473 X0.n941 X0.n254 2.2505
R17474 X0.n950 X0.n949 2.2505
R17475 X0.n252 X0.n249 2.2505
R17476 X0.n965 X0.n964 2.2505
R17477 X0.n963 X0.n962 2.2505
R17478 X0.n956 X0.n240 2.2505
R17479 X0.n978 X0.n235 2.2505
R17480 X0.n996 X0.n995 2.2505
R17481 X0.n984 X0.n233 2.2505
R17482 X0.n1001 X0.n1000 2.2505
R17483 X0.n1003 X0.n218 2.2505
R17484 X0.n1016 X0.n1015 2.2505
R17485 X0.n220 X0.n216 2.2505
R17486 X0.n1031 X0.n1030 2.2505
R17487 X0.n1029 X0.n1028 2.2505
R17488 X0.n1025 X0.n1022 2.2505
R17489 X0.n1042 X0.n200 2.2505
R17490 X0.n1057 X0.n1056 2.2505
R17491 X0.n1048 X0.n198 2.2505
R17492 X0.n1062 X0.n1061 2.2505
R17493 X0.n1065 X0.n187 2.2505
R17494 X0.n1083 X0.n1082 2.2505
R17495 X0.n1073 X0.n185 2.2505
R17496 X0.n1088 X0.n1087 2.2505
R17497 X0.n1091 X0.n173 2.2505
R17498 X0.n1114 X0.n1113 2.2505
R17499 X0.n1105 X0.n171 2.2505
R17500 X0.n1119 X0.n1118 2.2505
R17501 X0.n710 X0.n29 2.2505
R17502 X0.n1344 X0.n32 2.2505
R17503 X0.n1343 X0.n33 2.2505
R17504 X0.n1342 X0.n34 2.2505
R17505 X0.n693 X0.n35 2.2505
R17506 X0.n1338 X0.n37 2.2505
R17507 X0.n1337 X0.n38 2.2505
R17508 X0.n1336 X0.n39 2.2505
R17509 X0.n676 X0.n40 2.2505
R17510 X0.n1332 X0.n42 2.2505
R17511 X0.n1331 X0.n43 2.2505
R17512 X0.n1330 X0.n44 2.2505
R17513 X0.n538 X0.n45 2.2505
R17514 X0.n1326 X0.n47 2.2505
R17515 X0.n1325 X0.n48 2.2505
R17516 X0.n1324 X0.n49 2.2505
R17517 X0.n644 X0.n50 2.2505
R17518 X0.n1320 X0.n52 2.2505
R17519 X0.n1319 X0.n53 2.2505
R17520 X0.n1318 X0.n54 2.2505
R17521 X0.n629 X0.n55 2.2505
R17522 X0.n1314 X0.n57 2.2505
R17523 X0.n1313 X0.n58 2.2505
R17524 X0.n1312 X0.n59 2.2505
R17525 X0.n615 X0.n60 2.2505
R17526 X0.n1308 X0.n62 2.2505
R17527 X0.n1307 X0.n63 2.2505
R17528 X0.n1306 X0.n64 2.2505
R17529 X0.n571 X0.n65 2.2505
R17530 X0.n1302 X0.n67 2.2505
R17531 X0.n1301 X0.n68 2.2505
R17532 X0.n1300 X0.n69 2.2505
R17533 X0.n580 X0.n70 2.2505
R17534 X0.n1296 X0.n72 2.2505
R17535 X0.n1297 X0.n1296 2.2505
R17536 X0.n1298 X0.n70 2.2505
R17537 X0.n1300 X0.n1299 2.2505
R17538 X0.n1301 X0.n66 2.2505
R17539 X0.n1303 X0.n1302 2.2505
R17540 X0.n1304 X0.n65 2.2505
R17541 X0.n1306 X0.n1305 2.2505
R17542 X0.n1307 X0.n61 2.2505
R17543 X0.n1309 X0.n1308 2.2505
R17544 X0.n1310 X0.n60 2.2505
R17545 X0.n1312 X0.n1311 2.2505
R17546 X0.n1313 X0.n56 2.2505
R17547 X0.n1315 X0.n1314 2.2505
R17548 X0.n1316 X0.n55 2.2505
R17549 X0.n1318 X0.n1317 2.2505
R17550 X0.n1319 X0.n51 2.2505
R17551 X0.n1321 X0.n1320 2.2505
R17552 X0.n1322 X0.n50 2.2505
R17553 X0.n1324 X0.n1323 2.2505
R17554 X0.n1325 X0.n46 2.2505
R17555 X0.n1327 X0.n1326 2.2505
R17556 X0.n1328 X0.n45 2.2505
R17557 X0.n1330 X0.n1329 2.2505
R17558 X0.n1331 X0.n41 2.2505
R17559 X0.n1333 X0.n1332 2.2505
R17560 X0.n1334 X0.n40 2.2505
R17561 X0.n1336 X0.n1335 2.2505
R17562 X0.n1337 X0.n36 2.2505
R17563 X0.n1339 X0.n1338 2.2505
R17564 X0.n1340 X0.n35 2.2505
R17565 X0.n1342 X0.n1341 2.2505
R17566 X0.n1343 X0.n31 2.2505
R17567 X0.n1345 X0.n1344 2.2505
R17568 X0.n1346 X0.n29 2.2505
R17569 X0.n898 X0.n897 2.2505
R17570 X0.n895 X0.n894 2.2505
R17571 X0.n892 X0.n891 2.2505
R17572 X0.n889 X0.n888 2.2505
R17573 X0.n886 X0.n885 2.2505
R17574 X0.n1375 X0.n1374 2.2505
R17575 X0.n1372 X0.n1371 2.2505
R17576 X0.n1369 X0.n1368 2.2505
R17577 X0.n1367 X0.n11 2.2505
R17578 X0.n1364 X0.n15 2.2505
R17579 X0.n1361 X0.n16 2.2505
R17580 X0.n1358 X0.n20 2.2505
R17581 X0.n1355 X0.n21 2.2505
R17582 X0.n1352 X0.n25 2.2505
R17583 X0.n1349 X0.n26 2.2505
R17584 X0.n723 X0.n722 2.2005
R17585 X0.n728 X0.n512 2.2005
R17586 X0.n511 X0.n509 2.2005
R17587 X0.n736 X0.n735 2.2005
R17588 X0.n741 X0.n506 2.2005
R17589 X0.n505 X0.n503 2.2005
R17590 X0.n748 X0.n500 2.2005
R17591 X0.n499 X0.n497 2.2005
R17592 X0.n754 X0.n496 2.2005
R17593 X0.n495 X0.n493 2.2005
R17594 X0.n762 X0.n761 2.2005
R17595 X0.n767 X0.n490 2.2005
R17596 X0.n488 X0.n487 2.2005
R17597 X0.n774 X0.n486 2.2005
R17598 X0.n779 X0.n778 2.2005
R17599 X0.n781 X0.n780 2.2005
R17600 X0.n786 X0.n479 2.2005
R17601 X0.n478 X0.n476 2.2005
R17602 X0.n793 X0.n475 2.2005
R17603 X0.n799 X0.n798 2.2005
R17604 X0.n801 X0.n472 2.2005
R17605 X0.n806 X0.n805 2.2005
R17606 X0.n808 X0.n807 2.2005
R17607 X0.n814 X0.n813 2.2005
R17608 X0.n816 X0.n815 2.2005
R17609 X0.n821 X0.n458 2.2005
R17610 X0.n823 X0.n457 2.2005
R17611 X0.n828 X0.n454 2.2005
R17612 X0.n453 X0.n451 2.2005
R17613 X0.n835 X0.n446 2.2005
R17614 X0.n841 X0.n840 2.2005
R17615 X0.n844 X0.n843 2.2005
R17616 X0.n849 X0.n442 2.2005
R17617 X0.n851 X0.n441 2.2005
R17618 X0.n856 X0.n438 2.2005
R17619 X0.n437 X0.n435 2.2005
R17620 X0.n864 X0.n863 2.2005
R17621 X0.n869 X0.n432 2.2005
R17622 X0.n431 X0.n430 2.2005
R17623 X0.n876 X0.n427 2.2005
R17624 X0.n292 X0.n290 2.2005
R17625 X0.n883 X0.n882 2.2005
R17626 X0.n421 X0.n289 2.2005
R17627 X0.n415 X0.n414 2.2005
R17628 X0.n413 X0.n412 2.2005
R17629 X0.n407 X0.n406 2.2005
R17630 X0.n405 X0.n404 2.2005
R17631 X0.n400 X0.n399 2.2005
R17632 X0.n398 X0.n397 2.2005
R17633 X0.n391 X0.n390 2.2005
R17634 X0.n389 X0.n388 2.2005
R17635 X0.n381 X0.n380 2.2005
R17636 X0.n379 X0.n378 2.2005
R17637 X0.n372 X0.n371 2.2005
R17638 X0.n370 X0.n369 2.2005
R17639 X0.n364 X0.n363 2.2005
R17640 X0.n362 X0.n361 2.2005
R17641 X0.n355 X0.n317 2.2005
R17642 X0.n346 X0.n321 2.2005
R17643 X0.n348 X0.n347 2.2005
R17644 X0.n341 X0.n340 2.2005
R17645 X0.n75 X0.n74 2.2005
R17646 X0.n159 X0.n157 2.2005
R17647 X0.n1127 X0.n1126 2.2005
R17648 X0.n167 X0.n158 2.2005
R17649 X0.n166 X0.n165 2.2005
R17650 X0.n164 X0.n162 2.2005
R17651 X0.n160 X0.n153 2.2005
R17652 X0.n1135 X0.n152 2.2005
R17653 X0.n1139 X0.n1138 2.2005
R17654 X0.n1136 X0.n150 2.2005
R17655 X0.n1144 X0.n148 2.2005
R17656 X0.n1151 X0.n1150 2.2005
R17657 X0.n1149 X0.n149 2.2005
R17658 X0.n1147 X0.n1146 2.2005
R17659 X0.n143 X0.n142 2.2005
R17660 X0.n1164 X0.n1163 2.2005
R17661 X0.n1162 X0.n140 2.2005
R17662 X0.n1170 X0.n1169 2.2005
R17663 X0.n1171 X0.n138 2.2005
R17664 X0.n1173 X0.n1172 2.2005
R17665 X0.n1176 X0.n1175 2.2005
R17666 X0.n1177 X0.n136 2.2005
R17667 X0.n1180 X0.n1179 2.2005
R17668 X0.n134 X0.n131 2.2005
R17669 X0.n1189 X0.n1188 2.2005
R17670 X0.n1187 X0.n133 2.2005
R17671 X0.n1186 X0.n127 2.2005
R17672 X0.n1198 X0.n1197 2.2005
R17673 X0.n1199 X0.n125 2.2005
R17674 X0.n1202 X0.n1201 2.2005
R17675 X0.n1203 X0.n124 2.2005
R17676 X0.n1206 X0.n1205 2.2005
R17677 X0.n121 X0.n119 2.2005
R17678 X0.n1217 X0.n1216 2.2005
R17679 X0.n122 X0.n120 2.2005
R17680 X0.n1210 X0.n1209 2.2005
R17681 X0.n1211 X0.n114 2.2005
R17682 X0.n1226 X0.n113 2.2005
R17683 X0.n1228 X0.n1227 2.2005
R17684 X0.n1231 X0.n1230 2.2005
R17685 X0.n1232 X0.n110 2.2005
R17686 X0.n1235 X0.n1234 2.2005
R17687 X0.n111 X0.n105 2.2005
R17688 X0.n1250 X0.n1249 2.2005
R17689 X0.n1248 X0.n106 2.2005
R17690 X0.n1247 X0.n1246 2.2005
R17691 X0.n1244 X0.n1243 2.2005
R17692 X0.n1242 X0.n100 2.2005
R17693 X0.n1259 X0.n99 2.2005
R17694 X0.n1261 X0.n1260 2.2005
R17695 X0.n1264 X0.n1263 2.2005
R17696 X0.n1265 X0.n97 2.2005
R17697 X0.n1268 X0.n1267 2.2005
R17698 X0.n87 X0.n85 2.2005
R17699 X0.n1274 X0.n1273 2.2005
R17700 X0.n95 X0.n86 2.2005
R17701 X0.n94 X0.n93 2.2005
R17702 X0.n92 X0.n91 2.2005
R17703 X0.n90 X0.n81 2.2005
R17704 X0.n1283 X0.n80 2.2005
R17705 X0.n1286 X0.n1285 2.2005
R17706 X0.n327 X0.n277 2.2005
R17707 X0.n905 X0.n276 2.2005
R17708 X0.n907 X0.n906 2.2005
R17709 X0.n914 X0.n913 2.2005
R17710 X0.n915 X0.n270 2.2005
R17711 X0.n918 X0.n917 2.2005
R17712 X0.n920 X0.n268 2.2005
R17713 X0.n923 X0.n922 2.2005
R17714 X0.n264 X0.n263 2.2005
R17715 X0.n933 X0.n931 2.2005
R17716 X0.n259 X0.n258 2.2005
R17717 X0.n940 X0.n939 2.2005
R17718 X0.n943 X0.n942 2.2005
R17719 X0.n945 X0.n255 2.2005
R17720 X0.n948 X0.n947 2.2005
R17721 X0.n256 X0.n247 2.2005
R17722 X0.n968 X0.n967 2.2005
R17723 X0.n966 X0.n248 2.2005
R17724 X0.n251 X0.n250 2.2005
R17725 X0.n958 X0.n957 2.2005
R17726 X0.n961 X0.n960 2.2005
R17727 X0.n959 X0.n241 2.2005
R17728 X0.n976 X0.n975 2.2005
R17729 X0.n977 X0.n239 2.2005
R17730 X0.n980 X0.n979 2.2005
R17731 X0.n982 X0.n236 2.2005
R17732 X0.n994 X0.n993 2.2005
R17733 X0.n991 X0.n237 2.2005
R17734 X0.n986 X0.n985 2.2005
R17735 X0.n232 X0.n230 2.2005
R17736 X0.n1006 X0.n1005 2.2005
R17737 X0.n1004 X0.n231 2.2005
R17738 X0.n1002 X0.n227 2.2005
R17739 X0.n1011 X0.n219 2.2005
R17740 X0.n1014 X0.n1013 2.2005
R17741 X0.n222 X0.n221 2.2005
R17742 X0.n214 X0.n212 2.2005
R17743 X0.n1033 X0.n1032 2.2005
R17744 X0.n215 X0.n213 2.2005
R17745 X0.n1024 X0.n1023 2.2005
R17746 X0.n1027 X0.n1026 2.2005
R17747 X0.n207 X0.n205 2.2005
R17748 X0.n1041 X0.n1040 2.2005
R17749 X0.n1044 X0.n1043 2.2005
R17750 X0.n1046 X0.n201 2.2005
R17751 X0.n1055 X0.n1054 2.2005
R17752 X0.n1052 X0.n202 2.2005
R17753 X0.n1050 X0.n1049 2.2005
R17754 X0.n197 X0.n195 2.2005
R17755 X0.n1068 X0.n1067 2.2005
R17756 X0.n1066 X0.n196 2.2005
R17757 X0.n1064 X0.n1063 2.2005
R17758 X0.n191 X0.n188 2.2005
R17759 X0.n1081 X0.n1080 2.2005
R17760 X0.n1072 X0.n189 2.2005
R17761 X0.n1075 X0.n1074 2.2005
R17762 X0.n184 X0.n183 2.2005
R17763 X0.n1094 X0.n1093 2.2005
R17764 X0.n1092 X0.n181 2.2005
R17765 X0.n1090 X0.n1089 2.2005
R17766 X0.n178 X0.n174 2.2005
R17767 X0.n1112 X0.n1111 2.2005
R17768 X0.n177 X0.n175 2.2005
R17769 X0.n1107 X0.n1106 2.2005
R17770 X0.n1104 X0.n170 2.2005
R17771 X0.n709 X0.n523 2.2005
R17772 X0.n711 X0.n525 2.2005
R17773 X0.n713 X0.n712 2.2005
R17774 X0.n708 X0.n707 2.2005
R17775 X0.n706 X0.n705 2.2005
R17776 X0.n704 X0.n703 2.2005
R17777 X0.n702 X0.n701 2.2005
R17778 X0.n692 X0.n528 2.2005
R17779 X0.n694 X0.n531 2.2005
R17780 X0.n696 X0.n695 2.2005
R17781 X0.n691 X0.n690 2.2005
R17782 X0.n689 X0.n688 2.2005
R17783 X0.n687 X0.n686 2.2005
R17784 X0.n685 X0.n684 2.2005
R17785 X0.n674 X0.n533 2.2005
R17786 X0.n675 X0.n535 2.2005
R17787 X0.n679 X0.n678 2.2005
R17788 X0.n677 X0.n673 2.2005
R17789 X0.n671 X0.n670 2.2005
R17790 X0.n669 X0.n668 2.2005
R17791 X0.n667 X0.n666 2.2005
R17792 X0.n665 X0.n664 2.2005
R17793 X0.n663 X0.n662 2.2005
R17794 X0.n661 X0.n660 2.2005
R17795 X0.n659 X0.n658 2.2005
R17796 X0.n657 X0.n656 2.2005
R17797 X0.n655 X0.n654 2.2005
R17798 X0.n653 X0.n652 2.2005
R17799 X0.n545 X0.n540 2.2005
R17800 X0.n547 X0.n546 2.2005
R17801 X0.n647 X0.n646 2.2005
R17802 X0.n645 X0.n548 2.2005
R17803 X0.n643 X0.n642 2.2005
R17804 X0.n641 X0.n549 2.2005
R17805 X0.n640 X0.n639 2.2005
R17806 X0.n638 X0.n637 2.2005
R17807 X0.n636 X0.n635 2.2005
R17808 X0.n634 X0.n633 2.2005
R17809 X0.n632 X0.n631 2.2005
R17810 X0.n630 X0.n552 2.2005
R17811 X0.n628 X0.n627 2.2005
R17812 X0.n626 X0.n625 2.2005
R17813 X0.n624 X0.n623 2.2005
R17814 X0.n622 X0.n621 2.2005
R17815 X0.n620 X0.n619 2.2005
R17816 X0.n618 X0.n617 2.2005
R17817 X0.n616 X0.n556 2.2005
R17818 X0.n614 X0.n613 2.2005
R17819 X0.n612 X0.n557 2.2005
R17820 X0.n567 X0.n559 2.2005
R17821 X0.n569 X0.n568 2.2005
R17822 X0.n607 X0.n606 2.2005
R17823 X0.n605 X0.n604 2.2005
R17824 X0.n603 X0.n602 2.2005
R17825 X0.n601 X0.n600 2.2005
R17826 X0.n599 X0.n598 2.2005
R17827 X0.n597 X0.n596 2.2005
R17828 X0.n595 X0.n594 2.2005
R17829 X0.n593 X0.n592 2.2005
R17830 X0.n591 X0.n590 2.2005
R17831 X0.n589 X0.n588 2.2005
R17832 X0.n578 X0.n574 2.2005
R17833 X0.n579 X0.n577 2.2005
R17834 X0.n583 X0.n582 2.2005
R17835 X0.n581 X0.n76 2.2005
R17836 X0.n896 X0.n281 1.8005
R17837 X0.n310 X0.n283 1.8005
R17838 X0.n890 X0.n286 1.8005
R17839 X0.n297 X0.n288 1.8005
R17840 X0.n426 X0.n6 1.8005
R17841 X0.n1373 X0.n8 1.8005
R17842 X0.n842 X0.n10 1.8005
R17843 X0.n1366 X0.n14 1.8005
R17844 X0.n1362 X0.n17 1.8005
R17845 X0.n1360 X0.n19 1.8005
R17846 X0.n1356 X0.n22 1.8005
R17847 X0.n1354 X0.n24 1.8005
R17848 X0.n1350 X0.n27 1.8005
R17849 X0.n1282 X0.n1281 1.8005
R17850 X0.n1276 X0.n1275 1.8005
R17851 X0.n102 X0.n98 1.8005
R17852 X0.n1245 X0.n101 1.8005
R17853 X0.n1233 X0.n104 1.8005
R17854 X0.n1225 X0.n1224 1.8005
R17855 X0.n1204 X0.n118 1.8005
R17856 X0.n132 X0.n128 1.8005
R17857 X0.n1178 X0.n130 1.8005
R17858 X0.n145 X0.n139 1.8005
R17859 X0.n1145 X0.n144 1.8005
R17860 X0.n1137 X0.n147 1.8005
R17861 X0.n163 X0.n154 1.8005
R17862 X0.n1281 X0.n1280 1.8005
R17863 X0.n1277 X0.n1276 1.8005
R17864 X0.n1255 X0.n102 1.8005
R17865 X0.n1254 X0.n101 1.8005
R17866 X0.n104 X0.n103 1.8005
R17867 X0.n1224 X0.n1223 1.8005
R17868 X0.n118 X0.n117 1.8005
R17869 X0.n1193 X0.n128 1.8005
R17870 X0.n130 X0.n129 1.8005
R17871 X0.n1158 X0.n145 1.8005
R17872 X0.n1155 X0.n144 1.8005
R17873 X0.n147 X0.n146 1.8005
R17874 X0.n1131 X0.n154 1.8005
R17875 X0.n156 X0.n155 1.8005
R17876 X0.n1120 X0.n156 1.8005
R17877 X0.n1295 X0.n1294 1.8005
R17878 X0.n1295 X0.n71 1.8005
R17879 X0.n896 X0.n279 1.8005
R17880 X0.n893 X0.n283 1.8005
R17881 X0.n890 X0.n284 1.8005
R17882 X0.n887 X0.n288 1.8005
R17883 X0.n6 X0.n4 1.8005
R17884 X0.n1373 X0.n5 1.8005
R17885 X0.n1370 X0.n10 1.8005
R17886 X0.n1366 X0.n1365 1.8005
R17887 X0.n1363 X0.n1362 1.8005
R17888 X0.n1360 X0.n1359 1.8005
R17889 X0.n1357 X0.n1356 1.8005
R17890 X0.n1354 X0.n1353 1.8005
R17891 X0.n1351 X0.n1350 1.8005
R17892 X0.n899 X0.n278 1.5005
R17893 X0.n339 X0.n278 1.5005
R17894 X0.n1348 X0.n30 1.5005
R17895 X0.n1348 X0.n1347 1.5005
R17896 X0.n717 X0.n524 1.1125
R17897 X0.n1100 X0.n179 1.10836
R17898 X0.n1099 X0.n180 1.10443
R17899 X0.n1103 X0.n169 1.10381
R17900 X0.n719 X0.n718 1.10372
R17901 X0.n1095 X0.n182 1.10339
R17902 X0.n1111 X0.n1110 1.10272
R17903 X0.n1101 X0.n178 1.10272
R17904 X0.n1098 X0.n181 1.10272
R17905 X0.n716 X0.n525 1.10263
R17906 X0.n713 X0.n526 1.10263
R17907 X0.n1288 X0.n1287 1.1005
R17908 X0.n1125 X0.n1124 1.1005
R17909 X0.n161 X0.n151 1.1005
R17910 X0.n1141 X0.n1140 1.1005
R17911 X0.n1143 X0.n1142 1.1005
R17912 X0.n1148 X0.n141 1.1005
R17913 X0.n1166 X0.n1165 1.1005
R17914 X0.n1168 X0.n1167 1.1005
R17915 X0.n1174 X0.n135 1.1005
R17916 X0.n1182 X0.n1181 1.1005
R17917 X0.n1185 X0.n1184 1.1005
R17918 X0.n1183 X0.n126 1.1005
R17919 X0.n1200 X0.n123 1.1005
R17920 X0.n1207 X0.n1206 1.1005
R17921 X0.n1215 X0.n1214 1.1005
R17922 X0.n1213 X0.n1212 1.1005
R17923 X0.n1229 X0.n109 1.1005
R17924 X0.n1237 X0.n1236 1.1005
R17925 X0.n1238 X0.n107 1.1005
R17926 X0.n1239 X0.n108 1.1005
R17927 X0.n1241 X0.n1240 1.1005
R17928 X0.n1262 X0.n96 1.1005
R17929 X0.n1270 X0.n1269 1.1005
R17930 X0.n1272 X0.n1271 1.1005
R17931 X0.n88 X0.n79 1.1005
R17932 X0.n1123 X0.n1122 1.1005
R17933 X0.n908 X0.n274 1.1005
R17934 X0.n934 X0.n261 1.1005
R17935 X0.n989 X0.n988 1.1005
R17936 X0.n225 X0.n224 1.1005
R17937 X0.n1039 X0.n1038 1.1005
R17938 X0.n1109 X0.n1108 1.1005
R17939 X0.n1102 X0.n176 1.1005
R17940 X0.n1097 X0.n1096 1.1005
R17941 X0.n1077 X0.n1076 1.1005
R17942 X0.n1070 X0.n1069 1.1005
R17943 X0.n1037 X0.n206 1.1005
R17944 X0.n1035 X0.n1034 1.1005
R17945 X0.n226 X0.n211 1.1005
R17946 X0.n1008 X0.n1007 1.1005
R17947 X0.n990 X0.n229 1.1005
R17948 X0.n974 X0.n973 1.1005
R17949 X0.n970 X0.n969 1.1005
R17950 X0.n936 X0.n935 1.1005
R17951 X0.n912 X0.n911 1.1005
R17952 X0.n910 X0.n909 1.1005
R17953 X0.n336 X0.n329 1.1005
R17954 X0.n335 X0.n326 1.1005
R17955 X0.n328 X0.n275 1.1005
R17956 X0.n338 X0.n337 1.1005
R17957 X0.n724 X0.n723 1.1005
R17958 X0.n727 X0.n726 1.1005
R17959 X0.n728 X0.n510 1.1005
R17960 X0.n731 X0.n509 1.1005
R17961 X0.n734 X0.n508 1.1005
R17962 X0.n739 X0.n507 1.1005
R17963 X0.n741 X0.n740 1.1005
R17964 X0.n742 X0.n502 1.1005
R17965 X0.n747 X0.n746 1.1005
R17966 X0.n756 X0.n755 1.1005
R17967 X0.n757 X0.n493 1.1005
R17968 X0.n759 X0.n758 1.1005
R17969 X0.n765 X0.n491 1.1005
R17970 X0.n767 X0.n766 1.1005
R17971 X0.n768 X0.n489 1.1005
R17972 X0.n773 X0.n485 1.1005
R17973 X0.n784 X0.n480 1.1005
R17974 X0.n786 X0.n785 1.1005
R17975 X0.n787 X0.n477 1.1005
R17976 X0.n792 X0.n474 1.1005
R17977 X0.n794 X0.n793 1.1005
R17978 X0.n795 X0.n473 1.1005
R17979 X0.n800 X0.n471 1.1005
R17980 X0.n802 X0.n801 1.1005
R17981 X0.n805 X0.n804 1.1005
R17982 X0.n467 X0.n466 1.1005
R17983 X0.n811 X0.n464 1.1005
R17984 X0.n813 X0.n812 1.1005
R17985 X0.n465 X0.n463 1.1005
R17986 X0.n819 X0.n459 1.1005
R17987 X0.n827 X0.n826 1.1005
R17988 X0.n828 X0.n452 1.1005
R17989 X0.n831 X0.n451 1.1005
R17990 X0.n834 X0.n450 1.1005
R17991 X0.n838 X0.n448 1.1005
R17992 X0.n840 X0.n839 1.1005
R17993 X0.n449 X0.n447 1.1005
R17994 X0.n847 X0.n443 1.1005
R17995 X0.n855 X0.n854 1.1005
R17996 X0.n856 X0.n436 1.1005
R17997 X0.n859 X0.n435 1.1005
R17998 X0.n862 X0.n434 1.1005
R17999 X0.n867 X0.n433 1.1005
R18000 X0.n869 X0.n868 1.1005
R18001 X0.n870 X0.n429 1.1005
R18002 X0.n875 X0.n874 1.1005
R18003 X0.n423 X0.n422 1.1005
R18004 X0.n421 X0.n293 1.1005
R18005 X0.n420 X0.n419 1.1005
R18006 X0.n296 X0.n295 1.1005
R18007 X0.n412 X0.n411 1.1005
R18008 X0.n410 X0.n298 1.1005
R18009 X0.n300 X0.n299 1.1005
R18010 X0.n404 X0.n403 1.1005
R18011 X0.n401 X0.n400 1.1005
R18012 X0.n396 X0.n395 1.1005
R18013 X0.n393 X0.n392 1.1005
R18014 X0.n391 X0.n305 1.1005
R18015 X0.n385 X0.n306 1.1005
R18016 X0.n383 X0.n382 1.1005
R18017 X0.n381 X0.n308 1.1005
R18018 X0.n375 X0.n309 1.1005
R18019 X0.n374 X0.n311 1.1005
R18020 X0.n373 X0.n372 1.1005
R18021 X0.n369 X0.n368 1.1005
R18022 X0.n366 X0.n365 1.1005
R18023 X0.n359 X0.n319 1.1005
R18024 X0.n361 X0.n360 1.1005
R18025 X0.n358 X0.n318 1.1005
R18026 X0.n353 X0.n352 1.1005
R18027 X0.n343 X0.n323 1.1005
R18028 X0.n342 X0.n341 1.1005
R18029 X0.n333 X0.n332 1.1005
R18030 X0.n334 X0.n333 1.1005
R18031 X0.n331 X0.n326 1.1005
R18032 X0.n325 X0.n324 1.1005
R18033 X0.n351 X0.n321 1.1005
R18034 X0.n350 X0.n349 1.1005
R18035 X0.n348 X0.n322 1.1005
R18036 X0.n345 X0.n344 1.1005
R18037 X0.n354 X0.n320 1.1005
R18038 X0.n357 X0.n356 1.1005
R18039 X0.n316 X0.n315 1.1005
R18040 X0.n367 X0.n314 1.1005
R18041 X0.n313 X0.n312 1.1005
R18042 X0.n377 X0.n376 1.1005
R18043 X0.n384 X0.n307 1.1005
R18044 X0.n387 X0.n386 1.1005
R18045 X0.n394 X0.n304 1.1005
R18046 X0.n303 X0.n302 1.1005
R18047 X0.n402 X0.n301 1.1005
R18048 X0.n409 X0.n408 1.1005
R18049 X0.n417 X0.n416 1.1005
R18050 X0.n418 X0.n294 1.1005
R18051 X0.n424 X0.n291 1.1005
R18052 X0.n876 X0.n425 1.1005
R18053 X0.n878 X0.n877 1.1005
R18054 X0.n879 X0.n292 1.1005
R18055 X0.n881 X0.n880 1.1005
R18056 X0.n873 X0.n428 1.1005
R18057 X0.n872 X0.n871 1.1005
R18058 X0.n866 X0.n865 1.1005
R18059 X0.n861 X0.n860 1.1005
R18060 X0.n858 X0.n857 1.1005
R18061 X0.n849 X0.n848 1.1005
R18062 X0.n850 X0.n440 1.1005
R18063 X0.n852 X0.n851 1.1005
R18064 X0.n853 X0.n439 1.1005
R18065 X0.n846 X0.n845 1.1005
R18066 X0.n445 X0.n444 1.1005
R18067 X0.n837 X0.n836 1.1005
R18068 X0.n833 X0.n832 1.1005
R18069 X0.n830 X0.n829 1.1005
R18070 X0.n821 X0.n820 1.1005
R18071 X0.n822 X0.n456 1.1005
R18072 X0.n824 X0.n823 1.1005
R18073 X0.n825 X0.n455 1.1005
R18074 X0.n818 X0.n817 1.1005
R18075 X0.n461 X0.n460 1.1005
R18076 X0.n810 X0.n809 1.1005
R18077 X0.n470 X0.n468 1.1005
R18078 X0.n803 X0.n469 1.1005
R18079 X0.n797 X0.n796 1.1005
R18080 X0.n791 X0.n790 1.1005
R18081 X0.n789 X0.n788 1.1005
R18082 X0.n783 X0.n782 1.1005
R18083 X0.n775 X0.n774 1.1005
R18084 X0.n776 X0.n484 1.1005
R18085 X0.n778 X0.n777 1.1005
R18086 X0.n482 X0.n481 1.1005
R18087 X0.n772 X0.n771 1.1005
R18088 X0.n770 X0.n769 1.1005
R18089 X0.n764 X0.n763 1.1005
R18090 X0.n760 X0.n492 1.1005
R18091 X0.n754 X0.n494 1.1005
R18092 X0.n748 X0.n498 1.1005
R18093 X0.n750 X0.n749 1.1005
R18094 X0.n751 X0.n497 1.1005
R18095 X0.n753 X0.n752 1.1005
R18096 X0.n745 X0.n501 1.1005
R18097 X0.n744 X0.n743 1.1005
R18098 X0.n738 X0.n737 1.1005
R18099 X0.n733 X0.n732 1.1005
R18100 X0.n730 X0.n729 1.1005
R18101 X0.n725 X0.n513 1.1005
R18102 X0.n721 X0.n514 1.1005
R18103 X0.n521 X0.n515 1.1005
R18104 X0.n520 X0.n519 1.1005
R18105 X0.n1292 X0.n1291 1.1005
R18106 X0.n1290 X0.n78 1.1005
R18107 X0.n1289 X0.n78 1.1005
R18108 X0.n517 X0.n515 1.1005
R18109 X0.n519 X0.n518 1.1005
R18110 X0.n1293 X0.n77 1.1005
R18111 X0.n585 X0.n584 1.1005
R18112 X0.n587 X0.n586 1.1005
R18113 X0.n576 X0.n573 1.1005
R18114 X0.n575 X0.n572 1.1005
R18115 X0.n570 X0.n566 1.1005
R18116 X0.n609 X0.n608 1.1005
R18117 X0.n611 X0.n610 1.1005
R18118 X0.n565 X0.n558 1.1005
R18119 X0.n564 X0.n555 1.1005
R18120 X0.n563 X0.n554 1.1005
R18121 X0.n562 X0.n553 1.1005
R18122 X0.n561 X0.n551 1.1005
R18123 X0.n560 X0.n550 1.1005
R18124 X0.n642 X0.n544 1.1005
R18125 X0.n649 X0.n648 1.1005
R18126 X0.n651 X0.n650 1.1005
R18127 X0.n543 X0.n539 1.1005
R18128 X0.n542 X0.n537 1.1005
R18129 X0.n541 X0.n536 1.1005
R18130 X0.n672 X0.n534 1.1005
R18131 X0.n681 X0.n680 1.1005
R18132 X0.n683 X0.n682 1.1005
R18133 X0.n532 X0.n530 1.1005
R18134 X0.n698 X0.n697 1.1005
R18135 X0.n700 X0.n699 1.1005
R18136 X0.n529 X0.n527 1.1005
R18137 X0.n715 X0.n714 1.1005
R18138 X0.n720 X0.n522 1.1005
R18139 X0.n339 X0.n338 0.733833
R18140 X0.n1121 X0.n1120 0.733833
R18141 X0.n1294 X0.n1293 0.733833
R18142 X0.n720 X0.n30 0.733833
R18143 X0.n1038 X0.n204 0.573769
R18144 X0.n932 X0.n261 0.573769
R18145 X0.n224 X0.n223 0.573695
R18146 X0.n274 X0.n272 0.573695
R18147 X0.n988 X0.n987 0.573346
R18148 X0.n330 X0.n326 0.550549
R18149 X0.n516 X0.n515 0.550549
R18150 X0.n1037 X0.n208 0.39244
R18151 X0.n936 X0.n260 0.39244
R18152 X0.n1012 X0.n211 0.389994
R18153 X0.n910 X0.n273 0.389994
R18154 X0.n992 X0.n229 0.387191
R18155 X0.n1079 X0.n1078 0.384705
R18156 X0.n972 X0.n242 0.384705
R18157 X0.n1047 X0.n203 0.384705
R18158 X0.n937 X0.n257 0.384705
R18159 X0.n1071 X0.n193 0.382331
R18160 X0.n971 X0.n245 0.382331
R18161 X0.n1053 X0.n194 0.382034
R18162 X0.n944 X0.n246 0.382034
R18163 X0.n1036 X0.n209 0.379547
R18164 X0.n983 X0.n238 0.379547
R18165 X0.n919 X0.n262 0.379547
R18166 X0.n1010 X0.n1009 0.376968
R18167 X0.n1009 X0.n228 0.376876
R18168 X0.n1036 X0.n210 0.375976
R18169 X0.n921 X0.n262 0.375976
R18170 X0.n981 X0.n238 0.375884
R18171 X0.n1051 X0.n194 0.374982
R18172 X0.n946 X0.n246 0.374982
R18173 X0.n1071 X0.n192 0.374889
R18174 X0.n971 X0.n244 0.374889
R18175 X0.n1078 X0.n190 0.373984
R18176 X0.n972 X0.n243 0.373984
R18177 X0.n1045 X0.n203 0.373891
R18178 X0.n938 X0.n937 0.373891
R18179 X0.n1121 X0.n168 0.275034
R18180 X0 X0.n1376 0.253431
R18181 X0.n3 X0.n2 0.182739
R18182 X0.n2 X0 0.0563209
R18183 X0.n897 X0.n896 0.0405
R18184 X0.n896 X0.n895 0.0405
R18185 X0.n895 X0.n283 0.0405
R18186 X0.n891 X0.n283 0.0405
R18187 X0.n891 X0.n890 0.0405
R18188 X0.n890 X0.n889 0.0405
R18189 X0.n889 X0.n288 0.0405
R18190 X0.n885 X0.n288 0.0405
R18191 X0.n885 X0.n6 0.0405
R18192 X0.n1374 X0.n6 0.0405
R18193 X0.n1374 X0.n1373 0.0405
R18194 X0.n1373 X0.n1372 0.0405
R18195 X0.n1372 X0.n10 0.0405
R18196 X0.n1368 X0.n10 0.0405
R18197 X0.n1367 X0.n1366 0.0405
R18198 X0.n1366 X0.n15 0.0405
R18199 X0.n1362 X0.n15 0.0405
R18200 X0.n1362 X0.n1361 0.0405
R18201 X0.n1361 X0.n1360 0.0405
R18202 X0.n1360 X0.n20 0.0405
R18203 X0.n1356 X0.n20 0.0405
R18204 X0.n1356 X0.n1355 0.0405
R18205 X0.n1355 X0.n1354 0.0405
R18206 X0.n1354 X0.n25 0.0405
R18207 X0.n1350 X0.n25 0.0405
R18208 X0.n1350 X0.n1349 0.0405
R18209 X0.n1129 X0.n154 0.0405
R18210 X0.n1133 X0.n154 0.0405
R18211 X0.n1133 X0.n147 0.0405
R18212 X0.n1153 X0.n147 0.0405
R18213 X0.n1153 X0.n144 0.0405
R18214 X0.n1160 X0.n144 0.0405
R18215 X0.n1160 X0.n145 0.0405
R18216 X0.n1156 X0.n145 0.0405
R18217 X0.n1156 X0.n130 0.0405
R18218 X0.n1191 X0.n130 0.0405
R18219 X0.n1191 X0.n128 0.0405
R18220 X0.n1195 X0.n128 0.0405
R18221 X0.n1195 X0.n118 0.0405
R18222 X0.n1219 X0.n118 0.0405
R18223 X0.n1224 X0.n115 0.0405
R18224 X0.n1224 X0.n116 0.0405
R18225 X0.n116 X0.n104 0.0405
R18226 X0.n1252 X0.n104 0.0405
R18227 X0.n1252 X0.n101 0.0405
R18228 X0.n1257 X0.n101 0.0405
R18229 X0.n1257 X0.n102 0.0405
R18230 X0.n102 X0.n84 0.0405
R18231 X0.n1276 X0.n84 0.0405
R18232 X0.n1276 X0.n82 0.0405
R18233 X0.n1281 X0.n82 0.0405
R18234 X0.n1281 X0.n73 0.0405
R18235 X0.n1131 X0.n1130 0.0405
R18236 X0.n1132 X0.n1131 0.0405
R18237 X0.n1132 X0.n146 0.0405
R18238 X0.n1154 X0.n146 0.0405
R18239 X0.n1155 X0.n1154 0.0405
R18240 X0.n1159 X0.n1155 0.0405
R18241 X0.n1159 X0.n1158 0.0405
R18242 X0.n1158 X0.n1157 0.0405
R18243 X0.n1157 X0.n129 0.0405
R18244 X0.n1192 X0.n129 0.0405
R18245 X0.n1193 X0.n1192 0.0405
R18246 X0.n1194 X0.n1193 0.0405
R18247 X0.n1194 X0.n117 0.0405
R18248 X0.n1220 X0.n117 0.0405
R18249 X0.n1223 X0.n1221 0.0405
R18250 X0.n1223 X0.n1222 0.0405
R18251 X0.n1222 X0.n103 0.0405
R18252 X0.n1253 X0.n103 0.0405
R18253 X0.n1254 X0.n1253 0.0405
R18254 X0.n1256 X0.n1254 0.0405
R18255 X0.n1256 X0.n1255 0.0405
R18256 X0.n1255 X0.n83 0.0405
R18257 X0.n1277 X0.n83 0.0405
R18258 X0.n1278 X0.n1277 0.0405
R18259 X0.n1280 X0.n1278 0.0405
R18260 X0.n1280 X0.n1279 0.0405
R18261 X0.n898 X0.n279 0.0405
R18262 X0.n894 X0.n279 0.0405
R18263 X0.n894 X0.n893 0.0405
R18264 X0.n893 X0.n892 0.0405
R18265 X0.n892 X0.n284 0.0405
R18266 X0.n888 X0.n284 0.0405
R18267 X0.n888 X0.n887 0.0405
R18268 X0.n887 X0.n886 0.0405
R18269 X0.n886 X0.n4 0.0405
R18270 X0.n1375 X0.n5 0.0405
R18271 X0.n1371 X0.n5 0.0405
R18272 X0.n1371 X0.n1370 0.0405
R18273 X0.n1370 X0.n1369 0.0405
R18274 X0.n1365 X0.n11 0.0405
R18275 X0.n1365 X0.n1364 0.0405
R18276 X0.n1364 X0.n1363 0.0405
R18277 X0.n1363 X0.n16 0.0405
R18278 X0.n1359 X0.n16 0.0405
R18279 X0.n1359 X0.n1358 0.0405
R18280 X0.n1358 X0.n1357 0.0405
R18281 X0.n1357 X0.n21 0.0405
R18282 X0.n1353 X0.n21 0.0405
R18283 X0.n1353 X0.n1352 0.0405
R18284 X0.n1352 X0.n1351 0.0405
R18285 X0.n1351 X0.n26 0.0405
R18286 X0.n1368 X0.n1367 0.0360676
R18287 X0.n1219 X0.n115 0.0360676
R18288 X0.n1221 X0.n1220 0.0360676
R18289 X0.n901 X0.n900 0.0360676
R18290 X0.n901 X0.n266 0.0360676
R18291 X0.n926 X0.n266 0.0360676
R18292 X0.n927 X0.n926 0.0360676
R18293 X0.n928 X0.n927 0.0360676
R18294 X0.n928 X0.n253 0.0360676
R18295 X0.n951 X0.n253 0.0360676
R18296 X0.n952 X0.n951 0.0360676
R18297 X0.n953 X0.n952 0.0360676
R18298 X0.n954 X0.n953 0.0360676
R18299 X0.n955 X0.n954 0.0360676
R18300 X0.n955 X0.n234 0.0360676
R18301 X0.n997 X0.n234 0.0360676
R18302 X0.n998 X0.n997 0.0360676
R18303 X0.n999 X0.n998 0.0360676
R18304 X0.n999 X0.n217 0.0360676
R18305 X0.n1017 X0.n217 0.0360676
R18306 X0.n1018 X0.n1017 0.0360676
R18307 X0.n1019 X0.n1018 0.0360676
R18308 X0.n1020 X0.n1019 0.0360676
R18309 X0.n1021 X0.n1020 0.0360676
R18310 X0.n1021 X0.n199 0.0360676
R18311 X0.n1058 X0.n199 0.0360676
R18312 X0.n1059 X0.n1058 0.0360676
R18313 X0.n1060 X0.n1059 0.0360676
R18314 X0.n1060 X0.n186 0.0360676
R18315 X0.n1084 X0.n186 0.0360676
R18316 X0.n1085 X0.n1084 0.0360676
R18317 X0.n1086 X0.n1085 0.0360676
R18318 X0.n1086 X0.n172 0.0360676
R18319 X0.n1115 X0.n172 0.0360676
R18320 X0.n1116 X0.n1115 0.0360676
R18321 X0.n1117 X0.n1116 0.0360676
R18322 X0.n903 X0.n902 0.0360676
R18323 X0.n902 X0.n267 0.0360676
R18324 X0.n925 X0.n267 0.0360676
R18325 X0.n925 X0.n265 0.0360676
R18326 X0.n929 X0.n265 0.0360676
R18327 X0.n929 X0.n254 0.0360676
R18328 X0.n950 X0.n254 0.0360676
R18329 X0.n950 X0.n252 0.0360676
R18330 X0.n964 X0.n252 0.0360676
R18331 X0.n964 X0.n963 0.0360676
R18332 X0.n963 X0.n956 0.0360676
R18333 X0.n956 X0.n235 0.0360676
R18334 X0.n996 X0.n235 0.0360676
R18335 X0.n996 X0.n233 0.0360676
R18336 X0.n1000 X0.n233 0.0360676
R18337 X0.n1000 X0.n218 0.0360676
R18338 X0.n1016 X0.n218 0.0360676
R18339 X0.n1016 X0.n216 0.0360676
R18340 X0.n1030 X0.n216 0.0360676
R18341 X0.n1030 X0.n1029 0.0360676
R18342 X0.n1029 X0.n1022 0.0360676
R18343 X0.n1022 X0.n200 0.0360676
R18344 X0.n1057 X0.n200 0.0360676
R18345 X0.n1057 X0.n198 0.0360676
R18346 X0.n1061 X0.n198 0.0360676
R18347 X0.n1061 X0.n187 0.0360676
R18348 X0.n1083 X0.n187 0.0360676
R18349 X0.n1083 X0.n185 0.0360676
R18350 X0.n1087 X0.n185 0.0360676
R18351 X0.n1087 X0.n173 0.0360676
R18352 X0.n1114 X0.n173 0.0360676
R18353 X0.n1114 X0.n171 0.0360676
R18354 X0.n1118 X0.n171 0.0360676
R18355 X0.n1344 X0.n29 0.0360676
R18356 X0.n1344 X0.n1343 0.0360676
R18357 X0.n1343 X0.n1342 0.0360676
R18358 X0.n1342 X0.n35 0.0360676
R18359 X0.n1338 X0.n35 0.0360676
R18360 X0.n1338 X0.n1337 0.0360676
R18361 X0.n1337 X0.n1336 0.0360676
R18362 X0.n1336 X0.n40 0.0360676
R18363 X0.n1332 X0.n40 0.0360676
R18364 X0.n1332 X0.n1331 0.0360676
R18365 X0.n1331 X0.n1330 0.0360676
R18366 X0.n1330 X0.n45 0.0360676
R18367 X0.n1326 X0.n45 0.0360676
R18368 X0.n1326 X0.n1325 0.0360676
R18369 X0.n1325 X0.n1324 0.0360676
R18370 X0.n1324 X0.n50 0.0360676
R18371 X0.n1320 X0.n50 0.0360676
R18372 X0.n1320 X0.n1319 0.0360676
R18373 X0.n1319 X0.n1318 0.0360676
R18374 X0.n1318 X0.n55 0.0360676
R18375 X0.n1314 X0.n55 0.0360676
R18376 X0.n1314 X0.n1313 0.0360676
R18377 X0.n1313 X0.n1312 0.0360676
R18378 X0.n1312 X0.n60 0.0360676
R18379 X0.n1308 X0.n60 0.0360676
R18380 X0.n1308 X0.n1307 0.0360676
R18381 X0.n1307 X0.n1306 0.0360676
R18382 X0.n1306 X0.n65 0.0360676
R18383 X0.n1302 X0.n65 0.0360676
R18384 X0.n1302 X0.n1301 0.0360676
R18385 X0.n1301 X0.n1300 0.0360676
R18386 X0.n1300 X0.n70 0.0360676
R18387 X0.n1296 X0.n70 0.0360676
R18388 X0.n1346 X0.n1345 0.0360676
R18389 X0.n1345 X0.n31 0.0360676
R18390 X0.n1341 X0.n31 0.0360676
R18391 X0.n1341 X0.n1340 0.0360676
R18392 X0.n1340 X0.n1339 0.0360676
R18393 X0.n1339 X0.n36 0.0360676
R18394 X0.n1335 X0.n36 0.0360676
R18395 X0.n1335 X0.n1334 0.0360676
R18396 X0.n1334 X0.n1333 0.0360676
R18397 X0.n1333 X0.n41 0.0360676
R18398 X0.n1329 X0.n41 0.0360676
R18399 X0.n1329 X0.n1328 0.0360676
R18400 X0.n1328 X0.n1327 0.0360676
R18401 X0.n1327 X0.n46 0.0360676
R18402 X0.n1323 X0.n46 0.0360676
R18403 X0.n1323 X0.n1322 0.0360676
R18404 X0.n1322 X0.n1321 0.0360676
R18405 X0.n1321 X0.n51 0.0360676
R18406 X0.n1317 X0.n51 0.0360676
R18407 X0.n1317 X0.n1316 0.0360676
R18408 X0.n1316 X0.n1315 0.0360676
R18409 X0.n1315 X0.n56 0.0360676
R18410 X0.n1311 X0.n56 0.0360676
R18411 X0.n1311 X0.n1310 0.0360676
R18412 X0.n1310 X0.n1309 0.0360676
R18413 X0.n1309 X0.n61 0.0360676
R18414 X0.n1305 X0.n61 0.0360676
R18415 X0.n1305 X0.n1304 0.0360676
R18416 X0.n1304 X0.n1303 0.0360676
R18417 X0.n1303 X0.n66 0.0360676
R18418 X0.n1299 X0.n66 0.0360676
R18419 X0.n1299 X0.n1298 0.0360676
R18420 X0.n1298 X0.n1297 0.0360676
R18421 X0.n1369 X0.n11 0.0360676
R18422 X0.n1376 X0.n4 0.031527
R18423 X0.n897 X0.n278 0.0234189
R18424 X0.n1129 X0.n156 0.0234189
R18425 X0.n1130 X0.n155 0.0234189
R18426 X0.n899 X0.n898 0.0234189
R18427 X0.n1349 X0.n1348 0.0233108
R18428 X0.n1295 X0.n73 0.0233108
R18429 X0.n1279 X0.n71 0.0233108
R18430 X0.n1347 X0.n26 0.0233108
R18431 X0.n900 X0.n899 0.0227703
R18432 X0.n903 X0.n278 0.0227703
R18433 X0.n1348 X0.n29 0.0227703
R18434 X0.n1347 X0.n1346 0.0227703
R18435 X0.n363 X0.n362 0.0188784
R18436 X0.n371 X0.n370 0.0188784
R18437 X0.n380 X0.n379 0.0188784
R18438 X0.n390 X0.n389 0.0188784
R18439 X0.n399 X0.n398 0.0188784
R18440 X0.n414 X0.n289 0.0188784
R18441 X0.n883 X0.n290 0.0188784
R18442 X0.n430 X0.n427 0.0188784
R18443 X0.n863 X0.n432 0.0188784
R18444 X0.n438 X0.n437 0.0188784
R18445 X0.n442 X0.n441 0.0188784
R18446 X0.n841 X0.n446 0.0188784
R18447 X0.n454 X0.n453 0.0188784
R18448 X0.n458 X0.n457 0.0188784
R18449 X0.n815 X0.n814 0.0188784
R18450 X0.n807 X0.n806 0.0188784
R18451 X0.n798 X0.n472 0.0188784
R18452 X0.n478 X0.n475 0.0188784
R18453 X0.n487 X0.n486 0.0188784
R18454 X0.n761 X0.n490 0.0188784
R18455 X0.n496 X0.n495 0.0188784
R18456 X0.n500 X0.n499 0.0188784
R18457 X0.n506 X0.n505 0.0188784
R18458 X0.n164 X0.n153 0.0188784
R18459 X0.n1138 X0.n1135 0.0188784
R18460 X0.n1136 X0.n148 0.0188784
R18461 X0.n1151 X0.n149 0.0188784
R18462 X0.n1146 X0.n143 0.0188784
R18463 X0.n1172 X0.n1171 0.0188784
R18464 X0.n1177 X0.n1176 0.0188784
R18465 X0.n1179 X0.n131 0.0188784
R18466 X0.n1189 X0.n133 0.0188784
R18467 X0.n1197 X0.n127 0.0188784
R18468 X0.n1202 X0.n125 0.0188784
R18469 X0.n1205 X0.n119 0.0188784
R18470 X0.n1217 X0.n120 0.0188784
R18471 X0.n1209 X0.n114 0.0188784
R18472 X0.n1227 X0.n1226 0.0188784
R18473 X0.n1232 X0.n1231 0.0188784
R18474 X0.n1234 X0.n105 0.0188784
R18475 X0.n1250 X0.n106 0.0188784
R18476 X0.n1260 X0.n1259 0.0188784
R18477 X0.n1265 X0.n1264 0.0188784
R18478 X0.n1267 X0.n85 0.0188784
R18479 X0.n1274 X0.n86 0.0188784
R18480 X0.n93 X0.n92 0.0188784
R18481 X0.n339 X0.n277 0.0188784
R18482 X0.n906 X0.n905 0.0188784
R18483 X0.n915 X0.n914 0.0188784
R18484 X0.n917 X0.n268 0.0188784
R18485 X0.n1002 X0.n219 0.0188784
R18486 X0.n1014 X0.n221 0.0188784
R18487 X0.n1032 X0.n214 0.0188784
R18488 X0.n1024 X0.n215 0.0188784
R18489 X0.n709 X0.n30 0.0188784
R18490 X0.n712 X0.n711 0.0188784
R18491 X0.n707 X0.n706 0.0188784
R18492 X0.n703 X0.n702 0.0188784
R18493 X0.n643 X0.n549 0.0188784
R18494 X0.n639 X0.n638 0.0188784
R18495 X0.n635 X0.n634 0.0188784
R18496 X0.n631 X0.n630 0.0188784
R18497 X0.n347 X0.n346 0.0187703
R18498 X0.n362 X0.n317 0.0187703
R18499 X0.n406 X0.n405 0.0187703
R18500 X0.n414 X0.n413 0.0187703
R18501 X0.n843 X0.n442 0.0187703
R18502 X0.n479 X0.n478 0.0187703
R18503 X0.n780 X0.n779 0.0187703
R18504 X0.n735 X0.n506 0.0187703
R18505 X0.n512 X0.n511 0.0187703
R18506 X0.n1127 X0.n158 0.0187703
R18507 X0.n165 X0.n164 0.0187703
R18508 X0.n1163 X0.n1162 0.0187703
R18509 X0.n1171 X0.n1170 0.0187703
R18510 X0.n1203 X0.n1202 0.0187703
R18511 X0.n1246 X0.n106 0.0187703
R18512 X0.n1244 X0.n100 0.0187703
R18513 X0.n92 X0.n81 0.0187703
R18514 X0.n1285 X0.n1283 0.0187703
R18515 X0.n931 X0.n264 0.0187703
R18516 X0.n940 X0.n258 0.0187703
R18517 X0.n942 X0.n255 0.0187703
R18518 X0.n948 X0.n256 0.0187703
R18519 X0.n967 X0.n966 0.0187703
R18520 X0.n958 X0.n251 0.0187703
R18521 X0.n961 X0.n959 0.0187703
R18522 X0.n977 X0.n976 0.0187703
R18523 X0.n979 X0.n236 0.0187703
R18524 X0.n994 X0.n237 0.0187703
R18525 X0.n985 X0.n232 0.0187703
R18526 X0.n1005 X0.n1004 0.0187703
R18527 X0.n1041 X0.n205 0.0187703
R18528 X0.n1043 X0.n201 0.0187703
R18529 X0.n1055 X0.n202 0.0187703
R18530 X0.n1049 X0.n197 0.0187703
R18531 X0.n1067 X0.n1066 0.0187703
R18532 X0.n1064 X0.n188 0.0187703
R18533 X0.n1081 X0.n189 0.0187703
R18534 X0.n1074 X0.n184 0.0187703
R18535 X0.n1093 X0.n1092 0.0187703
R18536 X0.n1090 X0.n174 0.0187703
R18537 X0.n1112 X0.n175 0.0187703
R18538 X0.n1106 X0.n170 0.0187703
R18539 X0.n695 X0.n694 0.0187703
R18540 X0.n690 X0.n689 0.0187703
R18541 X0.n686 X0.n685 0.0187703
R18542 X0.n675 X0.n674 0.0187703
R18543 X0.n678 X0.n677 0.0187703
R18544 X0.n670 X0.n669 0.0187703
R18545 X0.n666 X0.n665 0.0187703
R18546 X0.n662 X0.n661 0.0187703
R18547 X0.n658 X0.n657 0.0187703
R18548 X0.n654 X0.n653 0.0187703
R18549 X0.n546 X0.n545 0.0187703
R18550 X0.n646 X0.n645 0.0187703
R18551 X0.n625 X0.n624 0.0187703
R18552 X0.n621 X0.n620 0.0187703
R18553 X0.n617 X0.n616 0.0187703
R18554 X0.n614 X0.n557 0.0187703
R18555 X0.n568 X0.n567 0.0187703
R18556 X0.n606 X0.n605 0.0187703
R18557 X0.n602 X0.n601 0.0187703
R18558 X0.n598 X0.n597 0.0187703
R18559 X0.n594 X0.n593 0.0187703
R18560 X0.n590 X0.n589 0.0187703
R18561 X0.n579 X0.n578 0.0187703
R18562 X0.n582 X0.n581 0.0187703
R18563 X0.n370 X0.n282 0.0185541
R18564 X0.n504 X0.n500 0.0185541
R18565 X0.n1135 X0.n1134 0.0185541
R18566 X0.n89 X0.n86 0.0185541
R18567 X0.n923 X0.n269 0.0184459
R18568 X0.n1027 X0.n1025 0.0184459
R18569 X0.n693 X0.n692 0.0184459
R18570 X0.n628 X0.n57 0.0184459
R18571 X0.n842 X0.n841 0.0182297
R18572 X0.n1205 X0.n1204 0.0182297
R18573 X0.n924 X0.n923 0.0181216
R18574 X0.n1028 X0.n1027 0.0181216
R18575 X0.n692 X0.n34 0.0181216
R18576 X0.n629 X0.n628 0.0181216
R18577 X0.n406 X0.n297 0.0175811
R18578 X0.n780 X0.n19 0.0175811
R18579 X0.n1162 X0.n139 0.0175811
R18580 X0.n1245 X0.n1244 0.0175811
R18581 X0.n931 X0.n930 0.0173649
R18582 X0.n1042 X0.n1041 0.0173649
R18583 X0.n695 X0.n37 0.0173649
R18584 X0.n624 X0.n58 0.0173649
R18585 X0.n917 X0.n916 0.0170405
R18586 X0.n1031 X0.n215 0.0170405
R18587 X0.n703 X0.n33 0.0170405
R18588 X0.n631 X0.n54 0.0170405
R18589 X0.n884 X0.n883 0.0167162
R18590 X0.n798 X0.n18 0.0167162
R18591 X0.n1176 X0.n137 0.0167162
R18592 X0.n1251 X0.n105 0.0167162
R18593 X0.n941 X0.n940 0.0162838
R18594 X0.n1056 X0.n201 0.0162838
R18595 X0.n689 X0.n38 0.0162838
R18596 X0.n620 X0.n59 0.0162838
R18597 X0.n438 X0.n9 0.0159595
R18598 X0.n457 X0.n13 0.0159595
R18599 X0.n1197 X0.n1196 0.0159595
R18600 X0.n1209 X0.n1208 0.0159595
R18601 X0.n914 X0.n271 0.0159595
R18602 X0.n220 X0.n214 0.0159595
R18603 X0.n707 X0.n32 0.0159595
R18604 X0.n635 X0.n53 0.0159595
R18605 X0.n346 X0.n281 0.0157432
R18606 X0.n511 X0.n27 0.0157432
R18607 X0.n163 X0.n158 0.0157432
R18608 X0.n1283 X0.n1282 0.0157432
R18609 X0.n379 X0.n310 0.0152027
R18610 X0.n496 X0.n24 0.0152027
R18611 X0.n1137 X0.n1136 0.0152027
R18612 X0.n1275 X0.n85 0.0152027
R18613 X0.n949 X0.n255 0.0152027
R18614 X0.n1048 X0.n202 0.0152027
R18615 X0.n685 X0.n39 0.0152027
R18616 X0.n616 X0.n615 0.0152027
R18617 X0.n453 X0.n12 0.0148784
R18618 X0.n1218 X0.n1217 0.0148784
R18619 X0.n905 X0.n904 0.0148784
R18620 X0.n1015 X0.n1014 0.0148784
R18621 X0.n711 X0.n710 0.0148784
R18622 X0.n639 X0.n52 0.0148784
R18623 X0.n399 X0.n287 0.0141216
R18624 X0.n486 X0.n483 0.0141216
R18625 X0.n1161 X0.n143 0.0141216
R18626 X0.n1259 X0.n1258 0.0141216
R18627 X0.n256 X0.n249 0.0141216
R18628 X0.n1062 X0.n197 0.0141216
R18629 X0.n676 X0.n675 0.0141216
R18630 X0.n557 X0.n62 0.0141216
R18631 X0.n1117 X0.n155 0.0137973
R18632 X0.n1118 X0.n156 0.0137973
R18633 X0.n1003 X0.n1002 0.0137973
R18634 X0.n1120 X0.n1119 0.0137973
R18635 X0.n644 X0.n643 0.0137973
R18636 X0.n1294 X0.n72 0.0137973
R18637 X0.n1296 X0.n1295 0.0137973
R18638 X0.n1297 X0.n71 0.0137973
R18639 X0.n585 X0.n77 0.0134381
R18640 X0.n427 X0.n426 0.0133649
R18641 X0.n806 X0.n17 0.0133649
R18642 X0.n1179 X0.n1178 0.0133649
R18643 X0.n1233 X0.n1232 0.0133649
R18644 X0.n966 X0.n965 0.0130405
R18645 X0.n1066 X0.n1065 0.0130405
R18646 X0.n677 X0.n42 0.0130405
R18647 X0.n568 X0.n63 0.0130405
R18648 X0.n1005 X0.n1001 0.0128243
R18649 X0.n1106 X0.n1105 0.0128243
R18650 X0.n646 X0.n49 0.0128243
R18651 X0.n582 X0.n580 0.0128243
R18652 X0.n863 X0.n8 0.0126081
R18653 X0.n815 X0.n14 0.0126081
R18654 X0.n133 X0.n132 0.0126081
R18655 X0.n1226 X0.n1225 0.0126081
R18656 X0.n340 X0.n280 0.0123919
R18657 X0.n722 X0.n28 0.0123919
R18658 X0.n1128 X0.n157 0.0123919
R18659 X0.n1284 X0.n74 0.0123919
R18660 X0.n962 X0.n958 0.0119595
R18661 X0.n1082 X0.n188 0.0119595
R18662 X0.n669 X0.n43 0.0119595
R18663 X0.n605 X0.n64 0.0119595
R18664 X0.n389 X0.n285 0.0118514
R18665 X0.n761 X0.n23 0.0118514
R18666 X0.n1152 X0.n1151 0.0118514
R18667 X0.n1266 X0.n1265 0.0118514
R18668 X0.n985 X0.n984 0.0117432
R18669 X0.n1113 X0.n1112 0.0117432
R18670 X0.n545 X0.n48 0.0117432
R18671 X0.n578 X0.n69 0.0117432
R18672 X0.n1123 X0.n168 0.0116588
R18673 X0.n340 X0.n339 0.011527
R18674 X0.n1120 X0.n157 0.011527
R18675 X0.n722 X0.n30 0.0114189
R18676 X0.n1294 X0.n74 0.0114189
R18677 X0.n699 X0.n529 0.0109762
R18678 X0.n698 X0.n530 0.0109762
R18679 X0.n682 X0.n681 0.0109762
R18680 X0.n541 X0.n534 0.0109762
R18681 X0.n543 X0.n542 0.0109762
R18682 X0.n650 X0.n649 0.0109762
R18683 X0.n560 X0.n544 0.0109762
R18684 X0.n562 X0.n561 0.0109762
R18685 X0.n564 X0.n563 0.0109762
R18686 X0.n610 X0.n565 0.0109762
R18687 X0.n609 X0.n566 0.0109762
R18688 X0.n576 X0.n575 0.0109762
R18689 X0.n586 X0.n585 0.0109762
R18690 X0.n1124 X0.n151 0.0109762
R18691 X0.n1141 X0.n151 0.0109762
R18692 X0.n1142 X0.n1141 0.0109762
R18693 X0.n1142 X0.n141 0.0109762
R18694 X0.n1166 X0.n141 0.0109762
R18695 X0.n1167 X0.n1166 0.0109762
R18696 X0.n1167 X0.n135 0.0109762
R18697 X0.n1182 X0.n135 0.0109762
R18698 X0.n1184 X0.n1182 0.0109762
R18699 X0.n1184 X0.n1183 0.0109762
R18700 X0.n1183 X0.n123 0.0109762
R18701 X0.n1214 X0.n1207 0.0109762
R18702 X0.n1214 X0.n1213 0.0109762
R18703 X0.n1213 X0.n109 0.0109762
R18704 X0.n1237 X0.n109 0.0109762
R18705 X0.n1238 X0.n1237 0.0109762
R18706 X0.n1239 X0.n1238 0.0109762
R18707 X0.n1240 X0.n1239 0.0109762
R18708 X0.n1240 X0.n96 0.0109762
R18709 X0.n1270 X0.n96 0.0109762
R18710 X0.n1271 X0.n1270 0.0109762
R18711 X0.n1271 X0.n79 0.0109762
R18712 X0.n1288 X0.n79 0.0109762
R18713 X0.n911 X0.n262 0.0109762
R18714 X0.n937 X0.n936 0.0109762
R18715 X0.n970 X0.n246 0.0109762
R18716 X0.n972 X0.n971 0.0109762
R18717 X0.n973 X0.n238 0.0109762
R18718 X0.n1008 X0.n229 0.0109762
R18719 X0.n1009 X0.n211 0.0109762
R18720 X0.n1036 X0.n1035 0.0109762
R18721 X0.n1037 X0.n203 0.0109762
R18722 X0.n1070 X0.n194 0.0109762
R18723 X0.n1078 X0.n1071 0.0109762
R18724 X0.n699 X0.n698 0.01095
R18725 X0.n682 X0.n530 0.01095
R18726 X0.n681 X0.n534 0.01095
R18727 X0.n542 X0.n541 0.01095
R18728 X0.n650 X0.n543 0.01095
R18729 X0.n649 X0.n544 0.01095
R18730 X0.n561 X0.n560 0.01095
R18731 X0.n563 X0.n562 0.01095
R18732 X0.n565 X0.n564 0.01095
R18733 X0.n610 X0.n609 0.01095
R18734 X0.n575 X0.n566 0.01095
R18735 X0.n586 X0.n576 0.01095
R18736 X0.n1207 X0.n123 0.01095
R18737 X0.n1289 X0.n1288 0.01095
R18738 X0.n911 X0.n910 0.01095
R18739 X0.n936 X0.n262 0.01095
R18740 X0.n937 X0.n246 0.01095
R18741 X0.n971 X0.n970 0.01095
R18742 X0.n973 X0.n972 0.01095
R18743 X0.n238 X0.n229 0.01095
R18744 X0.n1009 X0.n1008 0.01095
R18745 X0.n1035 X0.n211 0.01095
R18746 X0.n1037 X0.n1036 0.01095
R18747 X0.n203 X0.n194 0.01095
R18748 X0.n1071 X0.n1070 0.01095
R18749 X0.n1078 X0.n1077 0.01095
R18750 X0.n959 X0.n240 0.0108784
R18751 X0.n1073 X0.n189 0.0108784
R18752 X0.n665 X0.n44 0.0108784
R18753 X0.n601 X0.n571 0.0108784
R18754 X0.n390 X0.n286 0.0107703
R18755 X0.n490 X0.n22 0.0107703
R18756 X0.n1145 X0.n149 0.0107703
R18757 X0.n1264 X0.n98 0.0107703
R18758 X0.n995 X0.n994 0.0106622
R18759 X0.n1091 X0.n1090 0.0106622
R18760 X0.n654 X0.n47 0.0106622
R18761 X0.n590 X0.n68 0.0106622
R18762 X0.n1124 X0.n1123 0.0106095
R18763 X0.n432 X0.n7 0.0100135
R18764 X0.n814 X0.n462 0.0100135
R18765 X0.n1190 X0.n1189 0.0100135
R18766 X0.n1227 X0.n112 0.0100135
R18767 X0.n978 X0.n977 0.0097973
R18768 X0.n1088 X0.n184 0.0097973
R18769 X0.n661 X0.n538 0.0097973
R18770 X0.n597 X0.n67 0.0097973
R18771 X0.n1103 X0.n168 0.00967266
R18772 X0.n979 X0.n978 0.00958108
R18773 X0.n1093 X0.n1088 0.00958108
R18774 X0.n658 X0.n538 0.00958108
R18775 X0.n594 X0.n67 0.00958108
R18776 X0.n1376 X0.n1375 0.00947297
R18777 X0.n430 X0.n7 0.00925676
R18778 X0.n807 X0.n462 0.00925676
R18779 X0.n1190 X0.n131 0.00925676
R18780 X0.n1231 X0.n112 0.00925676
R18781 X0.n988 X0.n229 0.00880612
R18782 X0.n995 X0.n236 0.00871622
R18783 X0.n1092 X0.n1091 0.00871622
R18784 X0.n657 X0.n47 0.00871622
R18785 X0.n593 X0.n68 0.00871622
R18786 X0.n398 X0.n286 0.0085
R18787 X0.n487 X0.n22 0.0085
R18788 X0.n1146 X0.n1145 0.0085
R18789 X0.n1260 X0.n98 0.0085
R18790 X0.n976 X0.n240 0.0085
R18791 X0.n1074 X0.n1073 0.0085
R18792 X0.n662 X0.n44 0.0085
R18793 X0.n598 X0.n571 0.0085
R18794 X0.n529 X0.n526 0.00809524
R18795 X0.n1110 X0.n1109 0.00778095
R18796 X0.n984 X0.n237 0.00763514
R18797 X0.n1113 X0.n174 0.00763514
R18798 X0.n653 X0.n48 0.00763514
R18799 X0.n589 X0.n69 0.00763514
R18800 X0.n380 X0.n285 0.00741892
R18801 X0.n495 X0.n23 0.00741892
R18802 X0.n1152 X0.n148 0.00741892
R18803 X0.n1267 X0.n1266 0.00741892
R18804 X0.n962 X0.n961 0.00741892
R18805 X0.n1082 X0.n1081 0.00741892
R18806 X0.n666 X0.n43 0.00741892
R18807 X0.n602 X0.n64 0.00741892
R18808 X0.n1077 X0.n182 0.00725714
R18809 X0.n1109 X0.n1103 0.00707381
R18810 X0.n347 X0.n280 0.00698649
R18811 X0.n512 X0.n28 0.00698649
R18812 X0.n1128 X0.n1127 0.00698649
R18813 X0.n1285 X0.n1284 0.00698649
R18814 X0.n910 X0.n275 0.00696162
R18815 X0.n1291 X0.n1289 0.00691667
R18816 X0.n437 X0.n8 0.00666216
R18817 X0.n458 X0.n14 0.00666216
R18818 X0.n132 X0.n127 0.00666216
R18819 X0.n1225 X0.n114 0.00666216
R18820 X0.n1001 X0.n232 0.00655405
R18821 X0.n1105 X0.n175 0.00655405
R18822 X0.n546 X0.n49 0.00655405
R18823 X0.n580 X0.n579 0.00655405
R18824 X0.n965 X0.n251 0.00633784
R18825 X0.n1065 X0.n1064 0.00633784
R18826 X0.n670 X0.n42 0.00633784
R18827 X0.n606 X0.n63 0.00633784
R18828 X0.n426 X0.n290 0.00590541
R18829 X0.n472 X0.n17 0.00590541
R18830 X0.n1178 X0.n1177 0.00590541
R18831 X0.n1234 X0.n1233 0.00590541
R18832 X0.n224 X0.n211 0.00588776
R18833 X0.n910 X0.n274 0.00588776
R18834 X0.n1004 X0.n1003 0.00547297
R18835 X0.n1119 X0.n170 0.00547297
R18836 X0.n645 X0.n644 0.00547297
R18837 X0.n581 X0.n72 0.00547297
R18838 X0.n967 X0.n249 0.00525676
R18839 X0.n1067 X0.n1062 0.00525676
R18840 X0.n678 X0.n676 0.00525676
R18841 X0.n567 X0.n62 0.00525676
R18842 X0.n405 X0.n287 0.00514865
R18843 X0.n779 X0.n483 0.00514865
R18844 X0.n1163 X0.n1161 0.00514865
R18845 X0.n1258 X0.n100 0.00514865
R18846 X0.n1290 X0.n77 0.00440238
R18847 X0.n446 X0.n12 0.00439189
R18848 X0.n1218 X0.n119 0.00439189
R18849 X0.n904 X0.n277 0.00439189
R18850 X0.n1015 X0.n219 0.00439189
R18851 X0.n710 X0.n709 0.00439189
R18852 X0.n549 X0.n52 0.00439189
R18853 X0.n1126 X0.n159 0.00425921
R18854 X0.n167 X0.n166 0.00425921
R18855 X0.n1150 X0.n1149 0.00425921
R18856 X0.n1147 X0.n142 0.00425921
R18857 X0.n1173 X0.n138 0.00425921
R18858 X0.n1175 X0.n136 0.00425921
R18859 X0.n1180 X0.n134 0.00425921
R18860 X0.n1188 X0.n1187 0.00425921
R18861 X0.n1206 X0.n121 0.00425921
R18862 X0.n1228 X0.n113 0.00425921
R18863 X0.n1230 X0.n110 0.00425921
R18864 X0.n1235 X0.n111 0.00425921
R18865 X0.n1249 X0.n1248 0.00425921
R18866 X0.n1261 X0.n99 0.00425921
R18867 X0.n1263 X0.n97 0.00425921
R18868 X0.n90 X0.n80 0.00425921
R18869 X0.n1286 X0.n75 0.00425921
R18870 X0.n975 X0.n241 0.00425921
R18871 X0.n980 X0.n239 0.00425921
R18872 X0.n1075 X0.n1072 0.00425921
R18873 X0.n1094 X0.n183 0.00425921
R18874 X0.n704 X0.n701 0.00425921
R18875 X0.n531 X0.n528 0.00425921
R18876 X0.n696 X0.n691 0.00425921
R18877 X0.n688 X0.n687 0.00425921
R18878 X0.n668 X0.n667 0.00425921
R18879 X0.n664 X0.n663 0.00425921
R18880 X0.n660 X0.n659 0.00425921
R18881 X0.n656 X0.n655 0.00425921
R18882 X0.n642 X0.n641 0.00425921
R18883 X0.n632 X0.n552 0.00425921
R18884 X0.n627 X0.n626 0.00425921
R18885 X0.n623 X0.n622 0.00425921
R18886 X0.n619 X0.n618 0.00425921
R18887 X0.n604 X0.n603 0.00425921
R18888 X0.n600 X0.n599 0.00425921
R18889 X0.n596 X0.n595 0.00425921
R18890 X0.n592 X0.n591 0.00425921
R18891 X0.n1099 X0.n1098 0.00424524
R18892 X0.n166 X0.n162 0.0042371
R18893 X0.n160 X0.n152 0.0042371
R18894 X0.n1139 X0.n150 0.0042371
R18895 X0.n1150 X0.n1144 0.0042371
R18896 X0.n1164 X0.n140 0.0042371
R18897 X0.n1169 X0.n138 0.0042371
R18898 X0.n1187 X0.n1186 0.0042371
R18899 X0.n1199 X0.n1198 0.0042371
R18900 X0.n1201 X0.n124 0.0042371
R18901 X0.n1206 X0.n124 0.0042371
R18902 X0.n1216 X0.n121 0.0042371
R18903 X0.n1210 X0.n122 0.0042371
R18904 X0.n1211 X0.n113 0.0042371
R18905 X0.n1248 X0.n1247 0.0042371
R18906 X0.n1243 X0.n1242 0.0042371
R18907 X0.n1268 X0.n97 0.0042371
R18908 X0.n1273 X0.n87 0.0042371
R18909 X0.n95 X0.n94 0.0042371
R18910 X0.n91 X0.n90 0.0042371
R18911 X0.n918 X0.n270 0.0042371
R18912 X0.n947 X0.n247 0.0042371
R18913 X0.n968 X0.n248 0.0042371
R18914 X0.n1006 X0.n231 0.0042371
R18915 X0.n1033 X0.n213 0.0042371
R18916 X0.n1050 X0.n195 0.0042371
R18917 X0.n1068 X0.n196 0.0042371
R18918 X0.n1111 X0.n177 0.0042371
R18919 X0.n1107 X0.n1104 0.0042371
R18920 X0.n713 X0.n708 0.0042371
R18921 X0.n705 X0.n704 0.0042371
R18922 X0.n687 X0.n684 0.0042371
R18923 X0.n535 X0.n533 0.0042371
R18924 X0.n679 X0.n673 0.0042371
R18925 X0.n671 X0.n668 0.0042371
R18926 X0.n655 X0.n652 0.0042371
R18927 X0.n547 X0.n540 0.0042371
R18928 X0.n647 X0.n548 0.0042371
R18929 X0.n642 X0.n548 0.0042371
R18930 X0.n641 X0.n640 0.0042371
R18931 X0.n637 X0.n636 0.0042371
R18932 X0.n633 X0.n632 0.0042371
R18933 X0.n618 X0.n556 0.0042371
R18934 X0.n613 X0.n612 0.0042371
R18935 X0.n569 X0.n559 0.0042371
R18936 X0.n607 X0.n604 0.0042371
R18937 X0.n591 X0.n588 0.0042371
R18938 X0.n577 X0.n574 0.0042371
R18939 X0.n583 X0.n76 0.0042371
R18940 X0.n1293 X0.n76 0.0042371
R18941 X0.n718 X0.n522 0.00423273
R18942 X0.n335 X0.n334 0.00422178
R18943 X0.n521 X0.n520 0.00422178
R18944 X0.n1097 X0.n182 0.00421905
R18945 X0.n949 X0.n948 0.00417568
R18946 X0.n1049 X0.n1048 0.00417568
R18947 X0.n674 X0.n39 0.00417568
R18948 X0.n615 X0.n614 0.00417568
R18949 X0.n161 X0.n160 0.00410442
R18950 X0.n94 X0.n88 0.00410442
R18951 X0.n371 X0.n310 0.00406757
R18952 X0.n499 X0.n24 0.00406757
R18953 X0.n1138 X0.n1137 0.00406757
R18954 X0.n1275 X0.n1274 0.00406757
R18955 X0.n987 X0.n230 0.00402269
R18956 X0.n922 X0.n260 0.00398793
R18957 X0.n1026 X0.n208 0.00398793
R18958 X0.n700 X0.n528 0.00397174
R18959 X0.n659 X0.n539 0.00397174
R18960 X0.n627 X0.n553 0.00397174
R18961 X0.n595 X0.n573 0.00397174
R18962 X0.n1185 X0.n134 0.00394963
R18963 X0.n1230 X0.n1229 0.00394963
R18964 X0.n913 X0.n272 0.00394626
R18965 X0.n223 X0.n212 0.00394626
R18966 X0.n327 X0.n273 0.00393696
R18967 X0.n1012 X0.n1011 0.00393696
R18968 X0.n932 X0.n259 0.00390294
R18969 X0.n1044 X0.n204 0.00390294
R18970 X0.n993 X0.n992 0.00389381
R18971 X0.n943 X0.n257 0.00385851
R18972 X0.n957 X0.n242 0.00385851
R18973 X0.n1054 X0.n1047 0.00385851
R18974 X0.n1079 X0.n191 0.00385851
R18975 X0.n944 X0.n943 0.00380768
R18976 X0.n1054 X0.n1053 0.00380768
R18977 X0.n957 X0.n245 0.00380053
R18978 X0.n193 X0.n191 0.00380053
R18979 X0.n1148 X0.n1147 0.00379484
R18980 X0.n1262 X0.n1261 0.00379484
R18981 X0.n720 X0.n719 0.00379484
R18982 X0.n1121 X0.n169 0.00377273
R18983 X0.n919 X0.n918 0.0037725
R18984 X0.n993 X0.n983 0.0037725
R18985 X0.n213 X0.n209 0.0037725
R18986 X0.n1101 X0.n1100 0.00374762
R18987 X0.n1011 X0.n1010 0.00372958
R18988 X0.n683 X0.n533 0.0037285
R18989 X0.n613 X0.n558 0.0037285
R18990 X0.n231 X0.n228 0.00372177
R18991 X0.n673 X0.n672 0.00370639
R18992 X0.n608 X0.n569 0.00370639
R18993 X0.n1110 X0.n1102 0.00369524
R18994 X0.n1168 X0.n140 0.00366216
R18995 X0.n1243 X0.n108 0.00366216
R18996 X0.n181 X0.n180 0.00366216
R18997 X0.n1096 X0.n1095 0.00364005
R18998 X0.n317 X0.n281 0.00363514
R18999 X0.n735 X0.n27 0.00363514
R19000 X0.n165 X0.n163 0.00363514
R19001 X0.n1282 X0.n81 0.00363514
R19002 X0.n717 X0.n716 0.00359048
R19003 X0.n981 X0.n980 0.00358532
R19004 X0.n334 X0.n330 0.00357902
R19005 X0.n520 X0.n516 0.00357902
R19006 X0.n922 X0.n921 0.00357098
R19007 X0.n1026 X0.n210 0.00357098
R19008 X0.n1175 X0.n1174 0.00348526
R19009 X0.n111 X0.n107 0.00348526
R19010 X0.n947 X0.n946 0.003457
R19011 X0.n1051 X0.n1050 0.003457
R19012 X0.n248 X0.n244 0.00344926
R19013 X0.n196 X0.n192 0.00344926
R19014 X0.n691 X0.n532 0.00344103
R19015 X0.n664 X0.n536 0.00344103
R19016 X0.n622 X0.n555 0.00344103
R19017 X0.n600 X0.n570 0.00344103
R19018 X0.n960 X0.n243 0.00343273
R19019 X0.n1080 X0.n190 0.00343273
R19020 X0.n939 X0.n938 0.00341839
R19021 X0.n1046 X0.n1045 0.00341839
R19022 X0.n1038 X0.n1037 0.00341837
R19023 X0.n936 X0.n261 0.00341837
R19024 X0.n715 X0.n526 0.00335476
R19025 X0.n1143 X0.n150 0.00335258
R19026 X0.n1269 X0.n87 0.00335258
R19027 X0.n938 X0.n259 0.0033136
R19028 X0.n1045 X0.n1044 0.0033136
R19029 X0.n441 X0.n9 0.00331081
R19030 X0.n454 X0.n13 0.00331081
R19031 X0.n1196 X0.n125 0.00331081
R19032 X0.n1208 X0.n120 0.00331081
R19033 X0.n906 X0.n271 0.00331081
R19034 X0.n221 X0.n220 0.00331081
R19035 X0.n712 X0.n32 0.00331081
R19036 X0.n638 X0.n53 0.00331081
R19037 X0.n250 X0.n244 0.00330444
R19038 X0.n1063 X0.n192 0.00330444
R19039 X0.n243 X0.n241 0.0032992
R19040 X0.n1072 X0.n190 0.0032992
R19041 X0.n946 X0.n945 0.00329663
R19042 X0.n1052 X0.n1051 0.00329663
R19043 X0.n179 X0.n178 0.00324201
R19044 X0.n1198 X0.n126 0.00319779
R19045 X0.n1212 X0.n1210 0.00319779
R19046 X0.n1111 X0.n176 0.00319779
R19047 X0.n651 X0.n540 0.00319779
R19048 X0.n587 X0.n574 0.00319779
R19049 X0.n913 X0.n912 0.00317568
R19050 X0.n1034 X0.n212 0.00317568
R19051 X0.n708 X0.n527 0.00317568
R19052 X0.n636 X0.n551 0.00317568
R19053 X0.n921 X0.n920 0.00316007
R19054 X0.n1023 X0.n210 0.00316007
R19055 X0.n982 X0.n981 0.00314581
R19056 X0.n525 X0.n524 0.00310934
R19057 X0.n942 X0.n941 0.00309459
R19058 X0.n1056 X0.n1055 0.00309459
R19059 X0.n686 X0.n38 0.00309459
R19060 X0.n617 X0.n59 0.00309459
R19061 X0.n1126 X0.n1125 0.003043
R19062 X0.n1287 X0.n1286 0.003043
R19063 X0.n1010 X0.n227 0.00302306
R19064 X0.n228 X0.n227 0.00300884
R19065 X0.n376 X0.n374 0.0029881
R19066 X0.n409 X0.n299 0.0029881
R19067 X0.n880 X0.n424 0.0029881
R19068 X0.n796 X0.n471 0.0029881
R19069 X0.n983 X0.n982 0.00298054
R19070 X0.n920 X0.n919 0.00298054
R19071 X0.n1023 X0.n209 0.00298054
R19072 X0.n783 X0.n481 0.0029619
R19073 X0.n752 X0.n494 0.0029619
R19074 X0.n250 X0.n245 0.00293083
R19075 X0.n1063 X0.n193 0.00293083
R19076 X0.n945 X0.n944 0.0029237
R19077 X0.n1053 X0.n1052 0.0029237
R19078 X0.n1200 X0.n1199 0.00291032
R19079 X0.n1215 X0.n122 0.00291032
R19080 X0.n1007 X0.n230 0.00291032
R19081 X0.n1108 X0.n177 0.00291032
R19082 X0.n714 X0.n713 0.00291032
R19083 X0.n648 X0.n547 0.00291032
R19084 X0.n637 X0.n550 0.00291032
R19085 X0.n584 X0.n577 0.00291032
R19086 X0.n939 X0.n257 0.00289527
R19087 X0.n1047 X0.n1046 0.00289527
R19088 X0.n960 X0.n242 0.00289527
R19089 X0.n1080 X0.n1079 0.00289527
R19090 X0.n332 X0.n330 0.00287188
R19091 X0.n518 X0.n516 0.00284569
R19092 X0.n992 X0.n991 0.00283826
R19093 X0.n1291 X0.n1290 0.00283095
R19094 X0.n276 X0.n273 0.00279542
R19095 X0.n1013 X0.n1012 0.00279542
R19096 X0.n263 X0.n260 0.00276679
R19097 X0.n208 X0.n207 0.00276679
R19098 X0.n1140 X0.n1139 0.00275553
R19099 X0.n1273 X0.n1272 0.00275553
R19100 X0.n1122 X0.n159 0.00273342
R19101 X0.n1293 X0.n75 0.00273342
R19102 X0.n332 X0.n331 0.00272619
R19103 X0.n331 X0.n324 0.00272619
R19104 X0.n350 X0.n322 0.00272619
R19105 X0.n352 X0.n351 0.00272619
R19106 X0.n360 X0.n359 0.00272619
R19107 X0.n368 X0.n312 0.00272619
R19108 X0.n373 X0.n312 0.00272619
R19109 X0.n375 X0.n308 0.00272619
R19110 X0.n383 X0.n308 0.00272619
R19111 X0.n385 X0.n305 0.00272619
R19112 X0.n393 X0.n305 0.00272619
R19113 X0.n401 X0.n302 0.00272619
R19114 X0.n402 X0.n401 0.00272619
R19115 X0.n411 X0.n410 0.00272619
R19116 X0.n411 X0.n295 0.00272619
R19117 X0.n419 X0.n293 0.00272619
R19118 X0.n423 X0.n293 0.00272619
R19119 X0.n879 X0.n878 0.00272619
R19120 X0.n874 X0.n425 0.00272619
R19121 X0.n868 X0.n867 0.00272619
R19122 X0.n859 X0.n858 0.00272619
R19123 X0.n858 X0.n436 0.00272619
R19124 X0.n852 X0.n440 0.00272619
R19125 X0.n848 X0.n440 0.00272619
R19126 X0.n848 X0.n847 0.00272619
R19127 X0.n839 X0.n838 0.00272619
R19128 X0.n831 X0.n830 0.00272619
R19129 X0.n830 X0.n452 0.00272619
R19130 X0.n824 X0.n456 0.00272619
R19131 X0.n820 X0.n456 0.00272619
R19132 X0.n820 X0.n819 0.00272619
R19133 X0.n812 X0.n465 0.00272619
R19134 X0.n812 X0.n811 0.00272619
R19135 X0.n804 X0.n470 0.00272619
R19136 X0.n804 X0.n803 0.00272619
R19137 X0.n794 X0.n474 0.00272619
R19138 X0.n785 X0.n784 0.00272619
R19139 X0.n777 X0.n776 0.00272619
R19140 X0.n775 X0.n485 0.00272619
R19141 X0.n766 X0.n765 0.00272619
R19142 X0.n757 X0.n756 0.00272619
R19143 X0.n756 X0.n494 0.00272619
R19144 X0.n751 X0.n750 0.00272619
R19145 X0.n750 X0.n498 0.00272619
R19146 X0.n746 X0.n498 0.00272619
R19147 X0.n740 X0.n502 0.00272619
R19148 X0.n740 X0.n739 0.00272619
R19149 X0.n732 X0.n731 0.00272619
R19150 X0.n731 X0.n730 0.00272619
R19151 X0.n724 X0.n514 0.00272619
R19152 X0.n518 X0.n517 0.00272619
R19153 X0.n342 X0.n324 0.0027
R19154 X0.n351 X0.n350 0.0027
R19155 X0.n360 X0.n358 0.0027
R19156 X0.n368 X0.n367 0.0027
R19157 X0.n376 X0.n375 0.0027
R19158 X0.n403 X0.n402 0.0027
R19159 X0.n878 X0.n425 0.0027
R19160 X0.n868 X0.n429 0.0027
R19161 X0.n860 X0.n859 0.0027
R19162 X0.n839 X0.n449 0.0027
R19163 X0.n832 X0.n831 0.0027
R19164 X0.n803 X0.n802 0.0027
R19165 X0.n795 X0.n794 0.0027
R19166 X0.n785 X0.n477 0.0027
R19167 X0.n776 X0.n775 0.0027
R19168 X0.n766 X0.n489 0.0027
R19169 X0.n758 X0.n757 0.0027
R19170 X0.n730 X0.n510 0.0027
R19171 X0.n517 X0.n514 0.0027
R19172 X0.n403 X0.n299 0.00264762
R19173 X0.n777 X0.n481 0.00264762
R19174 X0.n697 X0.n696 0.00264496
R19175 X0.n623 X0.n554 0.00264496
R19176 X0.n975 X0.n974 0.00262285
R19177 X0.n1076 X0.n1075 0.00262285
R19178 X0.n663 X0.n537 0.00262285
R19179 X0.n599 X0.n572 0.00262285
R19180 X0.n424 X0.n423 0.00262143
R19181 X0.n796 X0.n795 0.00262143
R19182 X0.n1181 X0.n136 0.00260074
R19183 X0.n1236 X0.n1235 0.00260074
R19184 X0.n378 X0.n311 0.00257862
R19185 X0.n754 X0.n753 0.00257862
R19186 X0.n802 X0.n471 0.00256905
R19187 X0.n884 X0.n289 0.00255405
R19188 X0.n475 X0.n18 0.00255405
R19189 X0.n1172 X0.n137 0.00255405
R19190 X0.n1251 X0.n1250 0.00255405
R19191 X0.n880 X0.n879 0.00254286
R19192 X0.n784 X0.n783 0.00254286
R19193 X0.n882 X0.n881 0.0025344
R19194 X0.n410 X0.n409 0.00251667
R19195 X0.n800 X0.n799 0.00251228
R19196 X0.n337 X0.n336 0.0024936
R19197 X0.n374 X0.n373 0.00246429
R19198 X0.n752 X0.n751 0.00246429
R19199 X0.n1165 X0.n1164 0.00244595
R19200 X0.n1242 X0.n1241 0.00244595
R19201 X0.n394 X0.n393 0.0024381
R19202 X0.n770 X0.n489 0.0024381
R19203 X0.n407 X0.n300 0.00242383
R19204 X0.n781 X0.n482 0.00242383
R19205 X0.n718 X0.n717 0.00238571
R19206 X0.n1100 X0.n1099 0.00238571
R19207 X0.n357 X0.n320 0.00238571
R19208 X0.n366 X0.n315 0.00238571
R19209 X0.n386 X0.n384 0.00238571
R19210 X0.n395 X0.n394 0.00238571
R19211 X0.n418 X0.n417 0.00238571
R19212 X0.n873 X0.n872 0.00238571
R19213 X0.n866 X0.n434 0.00238571
R19214 X0.n846 X0.n444 0.00238571
R19215 X0.n837 X0.n450 0.00238571
R19216 X0.n826 X0.n452 0.00238571
R19217 X0.n818 X0.n460 0.00238571
R19218 X0.n810 X0.n466 0.00238571
R19219 X0.n790 X0.n789 0.00238571
R19220 X0.n771 X0.n770 0.00238571
R19221 X0.n764 X0.n492 0.00238571
R19222 X0.n745 X0.n744 0.00238571
R19223 X0.n738 X0.n508 0.00238571
R19224 X0.n349 X0.n348 0.00237961
R19225 X0.n353 X0.n321 0.00237961
R19226 X0.n361 X0.n319 0.00237961
R19227 X0.n369 X0.n313 0.00237961
R19228 X0.n372 X0.n313 0.00237961
R19229 X0.n381 X0.n309 0.00237961
R19230 X0.n382 X0.n381 0.00237961
R19231 X0.n391 X0.n306 0.00237961
R19232 X0.n392 X0.n391 0.00237961
R19233 X0.n400 X0.n303 0.00237961
R19234 X0.n400 X0.n301 0.00237961
R19235 X0.n412 X0.n298 0.00237961
R19236 X0.n412 X0.n296 0.00237961
R19237 X0.n421 X0.n420 0.00237961
R19238 X0.n422 X0.n421 0.00237961
R19239 X0.n877 X0.n292 0.00237961
R19240 X0.n876 X0.n875 0.00237961
R19241 X0.n869 X0.n433 0.00237961
R19242 X0.n857 X0.n435 0.00237961
R19243 X0.n857 X0.n856 0.00237961
R19244 X0.n851 X0.n850 0.00237961
R19245 X0.n850 X0.n849 0.00237961
R19246 X0.n849 X0.n443 0.00237961
R19247 X0.n840 X0.n448 0.00237961
R19248 X0.n829 X0.n451 0.00237961
R19249 X0.n829 X0.n828 0.00237961
R19250 X0.n823 X0.n822 0.00237961
R19251 X0.n822 X0.n821 0.00237961
R19252 X0.n821 X0.n459 0.00237961
R19253 X0.n813 X0.n463 0.00237961
R19254 X0.n813 X0.n464 0.00237961
R19255 X0.n805 X0.n468 0.00237961
R19256 X0.n805 X0.n469 0.00237961
R19257 X0.n793 X0.n792 0.00237961
R19258 X0.n786 X0.n480 0.00237961
R19259 X0.n778 X0.n484 0.00237961
R19260 X0.n774 X0.n773 0.00237961
R19261 X0.n767 X0.n491 0.00237961
R19262 X0.n755 X0.n493 0.00237961
R19263 X0.n755 X0.n754 0.00237961
R19264 X0.n749 X0.n497 0.00237961
R19265 X0.n749 X0.n748 0.00237961
R19266 X0.n748 X0.n747 0.00237961
R19267 X0.n742 X0.n741 0.00237961
R19268 X0.n741 X0.n507 0.00237961
R19269 X0.n733 X0.n509 0.00237961
R19270 X0.n729 X0.n509 0.00237961
R19271 X0.n723 X0.n721 0.00237961
R19272 X0.n338 X0.n329 0.00237961
R19273 X0.n908 X0.n907 0.00237961
R19274 X0.n969 X0.n247 0.00237961
R19275 X0.n969 X0.n968 0.00237961
R19276 X0.n989 X0.n986 0.00237961
R19277 X0.n225 X0.n222 0.00237961
R19278 X0.n1069 X0.n195 0.00237961
R19279 X0.n1069 X0.n1068 0.00237961
R19280 X0.n680 X0.n535 0.00237961
R19281 X0.n680 X0.n679 0.00237961
R19282 X0.n612 X0.n611 0.00237961
R19283 X0.n611 X0.n559 0.00237961
R19284 X0.n872 X0.n429 0.00235952
R19285 X0.n853 X0.n852 0.00235952
R19286 X0.n341 X0.n325 0.00235749
R19287 X0.n349 X0.n321 0.00235749
R19288 X0.n361 X0.n318 0.00235749
R19289 X0.n369 X0.n314 0.00235749
R19290 X0.n377 X0.n309 0.00235749
R19291 X0.n404 X0.n301 0.00235749
R19292 X0.n877 X0.n876 0.00235749
R19293 X0.n870 X0.n869 0.00235749
R19294 X0.n861 X0.n435 0.00235749
R19295 X0.n840 X0.n447 0.00235749
R19296 X0.n833 X0.n451 0.00235749
R19297 X0.n801 X0.n469 0.00235749
R19298 X0.n793 X0.n473 0.00235749
R19299 X0.n787 X0.n786 0.00235749
R19300 X0.n774 X0.n484 0.00235749
R19301 X0.n768 X0.n767 0.00235749
R19302 X0.n759 X0.n493 0.00235749
R19303 X0.n729 X0.n728 0.00235749
R19304 X0.n934 X0.n933 0.00235749
R19305 X0.n1040 X0.n1039 0.00235749
R19306 X0.n811 X0.n810 0.00233333
R19307 X0.n404 X0.n300 0.00231327
R19308 X0.n778 X0.n482 0.00231327
R19309 X0.n343 X0.n342 0.00230714
R19310 X0.n726 X0.n510 0.00230714
R19311 X0.n725 X0.n724 0.00230714
R19312 X0.n422 X0.n291 0.00229115
R19313 X0.n797 X0.n473 0.00229115
R19314 X0.n1165 X0.n142 0.00229115
R19315 X0.n1241 X0.n99 0.00229115
R19316 X0.n344 X0.n322 0.00228095
R19317 X0.n359 X0.n315 0.00228095
R19318 X0.n744 X0.n502 0.00225476
R19319 X0.n801 X0.n800 0.00224693
R19320 X0.n916 X0.n915 0.00222973
R19321 X0.n1032 X0.n1031 0.00222973
R19322 X0.n706 X0.n33 0.00222973
R19323 X0.n634 X0.n54 0.00222973
R19324 X0.n881 X0.n292 0.00222482
R19325 X0.n782 X0.n480 0.00222482
R19326 X0.n408 X0.n298 0.0022027
R19327 X0.n854 X0.n436 0.00220238
R19328 X0.n825 X0.n824 0.00220238
R19329 X0.n449 X0.n444 0.00217619
R19330 X0.n838 X0.n837 0.00217619
R19331 X0.n372 X0.n311 0.00215848
R19332 X0.n753 X0.n497 0.00215848
R19333 X0.n392 X0.n304 0.00213636
R19334 X0.n769 X0.n768 0.00213636
R19335 X0.n1181 X0.n1180 0.00213636
R19336 X0.n1236 X0.n110 0.00213636
R19337 X0.n974 X0.n239 0.00211425
R19338 X0.n1076 X0.n183 0.00211425
R19339 X0.n660 X0.n537 0.00211425
R19340 X0.n596 X0.n572 0.00211425
R19341 X0.n716 X0.n715 0.00209762
R19342 X0.n358 X0.n357 0.00209762
R19343 X0.n828 X0.n827 0.00209214
R19344 X0.n935 X0.n263 0.00209214
R19345 X0.n207 X0.n206 0.00209214
R19346 X0.n697 X0.n531 0.00209214
R19347 X0.n626 X0.n554 0.00209214
R19348 X0.n739 X0.n738 0.00207143
R19349 X0.n871 X0.n870 0.00207002
R19350 X0.n851 X0.n439 0.00207002
R19351 X0.n809 X0.n464 0.00204791
R19352 X0.n341 X0.n323 0.0020258
R19353 X0.n728 X0.n727 0.0020258
R19354 X0.n723 X0.n513 0.0020258
R19355 X0.n867 X0.n866 0.00201905
R19356 X0.n930 X0.n258 0.00201351
R19357 X0.n1043 X0.n1042 0.00201351
R19358 X0.n690 X0.n37 0.00201351
R19359 X0.n621 X0.n58 0.00201351
R19360 X0.n348 X0.n345 0.00200369
R19361 X0.n319 X0.n316 0.00200369
R19362 X0.n1140 X0.n152 0.00200369
R19363 X0.n1272 X0.n95 0.00200369
R19364 X0.n337 X0.n335 0.00200107
R19365 X0.n336 X0.n275 0.00200107
R19366 X0.n522 X0.n521 0.00200107
R19367 X0.n465 X0.n460 0.00199286
R19368 X0.n743 X0.n742 0.00198157
R19369 X0.n856 X0.n855 0.00193735
R19370 X0.n823 X0.n455 0.00193735
R19371 X0.n447 X0.n445 0.00191523
R19372 X0.n836 X0.n448 0.00191523
R19373 X0.n338 X0.n326 0.00191523
R19374 X0.n329 X0.n328 0.00191523
R19375 X0.n720 X0.n515 0.00191523
R19376 X0.n1293 X0.n1292 0.00191523
R19377 X0.n386 X0.n385 0.00191429
R19378 X0.n765 X0.n764 0.00191429
R19379 X0.n397 X0.n396 0.00187101
R19380 X0.n933 X0.n932 0.00185493
R19381 X0.n1040 X0.n204 0.00185493
R19382 X0.n356 X0.n318 0.00184889
R19383 X0.n772 X0.n488 0.00184889
R19384 X0.n1201 X0.n1200 0.00184889
R19385 X0.n1216 X0.n1215 0.00184889
R19386 X0.n909 X0.n276 0.00184889
R19387 X0.n1007 X0.n1006 0.00184889
R19388 X0.n1013 X0.n226 0.00184889
R19389 X0.n1108 X0.n1107 0.00184889
R19390 X0.n714 X0.n525 0.00184889
R19391 X0.n648 X0.n647 0.00184889
R19392 X0.n640 X0.n550 0.00184889
R19393 X0.n584 X0.n583 0.00184889
R19394 X0.n789 X0.n477 0.00183571
R19395 X0.n737 X0.n507 0.00182678
R19396 X0.n417 X0.n295 0.00180952
R19397 X0.n413 X0.n297 0.0017973
R19398 X0.n479 X0.n19 0.0017973
R19399 X0.n1170 X0.n139 0.0017973
R19400 X0.n1246 X0.n1245 0.0017973
R19401 X0.n907 X0.n272 0.0017897
R19402 X0.n223 X0.n222 0.0017897
R19403 X0.n431 X0.n428 0.00178256
R19404 X0.n865 X0.n433 0.00178256
R19405 X0.n808 X0.n467 0.00178256
R19406 X0.n463 X0.n461 0.00176044
R19407 X0.n1102 X0.n1101 0.00175714
R19408 X0.n419 X0.n418 0.00173095
R19409 X0.n790 X0.n474 0.00173095
R19410 X0.n365 X0.n364 0.00171622
R19411 X0.n987 X0.n986 0.00171347
R19412 X0.n387 X0.n306 0.0016941
R19413 X0.n763 X0.n491 0.0016941
R19414 X0.n503 X0.n501 0.0016941
R19415 X0.n1125 X0.n167 0.0016941
R19416 X0.n1287 X0.n80 0.0016941
R19417 X0.n758 X0.n492 0.00165238
R19418 X0.n845 X0.n844 0.00162776
R19419 X0.n835 X0.n834 0.00162776
R19420 X0.n788 X0.n787 0.00162776
R19421 X0.n524 X0.n523 0.00162776
R19422 X0.n384 X0.n383 0.00162619
R19423 X0.n416 X0.n296 0.00160565
R19424 X0.n912 X0.n270 0.00158354
R19425 X0.n1034 X0.n1033 0.00158354
R19426 X0.n705 X0.n527 0.00158354
R19427 X0.n633 X0.n551 0.00158354
R19428 X0.n355 X0.n354 0.00156143
R19429 X0.n736 X0.n734 0.00156143
R19430 X0.n1186 X0.n126 0.00156143
R19431 X0.n1212 X0.n1211 0.00156143
R19432 X0.n991 X0.n990 0.00156143
R19433 X0.n178 X0.n176 0.00156143
R19434 X0.n652 X0.n651 0.00156143
R19435 X0.n588 X0.n587 0.00156143
R19436 X0.n860 X0.n434 0.00154762
R19437 X0.n819 X0.n818 0.00154762
R19438 X0.n420 X0.n294 0.00153931
R19439 X0.n792 X0.n791 0.00153931
R19440 X0.n864 X0.n862 0.00149509
R19441 X0.n1089 X0.n179 0.00149509
R19442 X0.n817 X0.n816 0.00147297
R19443 X0.n760 X0.n759 0.00147297
R19444 X0.n352 X0.n320 0.00146905
R19445 X0.n732 X0.n508 0.00146905
R19446 X0.n382 X0.n307 0.00145086
R19447 X0.n388 X0.n307 0.00140663
R19448 X0.n762 X0.n760 0.00140663
R19449 X0.n1144 X0.n1143 0.00140663
R19450 X0.n1269 X0.n1268 0.00140663
R19451 X0.n832 X0.n450 0.00139048
R19452 X0.n862 X0.n861 0.00138452
R19453 X0.n817 X0.n459 0.00138452
R19454 X0.n344 X0.n343 0.00136429
R19455 X0.n854 X0.n853 0.00136429
R19456 X0.n847 X0.n846 0.00136429
R19457 X0.n415 X0.n294 0.00134029
R19458 X0.n791 X0.n476 0.00134029
R19459 X0.n826 X0.n825 0.00133809
R19460 X0.n726 X0.n725 0.00133809
R19461 X0.n354 X0.n353 0.00131818
R19462 X0.n734 X0.n733 0.00131818
R19463 X0.n990 X0.n989 0.00131818
R19464 X0.n688 X0.n532 0.00129607
R19465 X0.n667 X0.n536 0.00129607
R19466 X0.n619 X0.n555 0.00129607
R19467 X0.n603 X0.n570 0.00129607
R19468 X0.n367 X0.n366 0.00128571
R19469 X0.n746 X0.n745 0.00128571
R19470 X0.n416 X0.n415 0.00125184
R19471 X0.n834 X0.n833 0.00125184
R19472 X0.n788 X0.n476 0.00125184
R19473 X0.n1174 X0.n1173 0.00125184
R19474 X0.n1249 X0.n107 0.00125184
R19475 X0.n345 X0.n323 0.00122973
R19476 X0.n855 X0.n439 0.00122973
R19477 X0.n845 X0.n443 0.00122973
R19478 X0.n827 X0.n455 0.00120762
R19479 X0.n727 X0.n513 0.00120762
R19480 X0.n874 X0.n873 0.00120714
R19481 X0.n470 X0.n466 0.00120714
R19482 X0.n388 X0.n387 0.0011855
R19483 X0.n763 X0.n762 0.0011855
R19484 X0.n365 X0.n314 0.00116339
R19485 X0.n747 X0.n501 0.00116339
R19486 X0.n924 X0.n268 0.00114865
R19487 X0.n1028 X0.n1024 0.00114865
R19488 X0.n702 X0.n34 0.00114865
R19489 X0.n630 X0.n629 0.00114865
R19490 X0.n771 X0.n485 0.00112857
R19491 X0.n816 X0.n461 0.00111916
R19492 X0.n395 X0.n302 0.00110238
R19493 X0.n875 X0.n428 0.00109705
R19494 X0.n865 X0.n864 0.00109705
R19495 X0.n468 X0.n467 0.00109705
R19496 X0.n1169 X0.n1168 0.00109705
R19497 X0.n1247 X0.n108 0.00109705
R19498 X0.n1089 X0.n180 0.00109705
R19499 X0.n672 X0.n671 0.00105283
R19500 X0.n608 X0.n607 0.00105283
R19501 X0.n1292 X0.n78 0.00105283
R19502 X0.n843 X0.n842 0.00104054
R19503 X0.n1204 X0.n1203 0.00104054
R19504 X0.n356 X0.n355 0.00103071
R19505 X0.n773 X0.n772 0.00103071
R19506 X0.n737 X0.n736 0.00103071
R19507 X0.n333 X0.n326 0.00103071
R19508 X0.n909 X0.n908 0.00103071
R19509 X0.n226 X0.n225 0.00103071
R19510 X0.n519 X0.n515 0.00103071
R19511 X0.n684 X0.n683 0.00103071
R19512 X0.n558 X0.n556 0.00103071
R19513 X0.n396 X0.n303 0.0010086
R19514 X0.n844 X0.n445 0.000964373
R19515 X0.n836 X0.n835 0.000964373
R19516 X0.n328 X0.n327 0.000964373
R19517 X0.n1104 X0.n169 0.000964373
R19518 X0.n719 X0.n523 0.000964373
R19519 X0.n1149 X0.n1148 0.00094226
R19520 X0.n1263 X0.n1262 0.00094226
R19521 X0.n269 X0.n264 0.000932432
R19522 X0.n1025 X0.n205 0.000932432
R19523 X0.n694 X0.n693 0.000932432
R19524 X0.n625 X0.n57 0.000932432
R19525 X0.n338 X0.n325 0.000898034
R19526 X0.n743 X0.n503 0.000898034
R19527 X0.n364 X0.n316 0.000875921
R19528 X0.n721 X0.n720 0.000853808
R19529 X0.n1095 X0.n1094 0.000831695
R19530 X0.n1098 X0.n1097 0.000814286
R19531 X0.n871 X0.n431 0.000809582
R19532 X0.n809 X0.n808 0.000809582
R19533 X0.n1188 X0.n1185 0.000787469
R19534 X0.n1229 X0.n1228 0.000787469
R19535 X0.n935 X0.n934 0.000787469
R19536 X0.n1039 X0.n206 0.000787469
R19537 X0.n1096 X0.n181 0.000765356
R19538 X0.n701 X0.n700 0.000765356
R19539 X0.n656 X0.n539 0.000765356
R19540 X0.n553 X0.n552 0.000765356
R19541 X0.n592 X0.n573 0.000765356
R19542 X0.n769 X0.n488 0.000743243
R19543 X0.n397 X0.n304 0.00072113
R19544 X0.n363 X0.n282 0.000716216
R19545 X0.n505 X0.n504 0.000716216
R19546 X0.n1134 X0.n153 0.000716216
R19547 X0.n93 X0.n89 0.000716216
R19548 X0.n408 X0.n407 0.000676904
R19549 X0.n782 X0.n781 0.000654791
R19550 X0.n162 X0.n161 0.000654791
R19551 X0.n91 X0.n88 0.000654791
R19552 X0.n799 X0.n797 0.000588452
R19553 X0.n882 X0.n291 0.000566339
R19554 X0.n378 X0.n377 0.000522113
R19555 X0.n1122 X0.n1121 0.000522113
R19556 VSS.n1142 VSS.n1141 1.1469e+07
R19557 VSS.n1108 VSS.n9 7.365e+06
R19558 VSS.n871 VSS.n870 6.74962e+06
R19559 VSS.n441 VSS.n9 6.543e+06
R19560 VSS.n9 VSS.n8 6.2235e+06
R19561 VSS.n1142 VSS.n416 5.286e+06
R19562 VSS.n1141 VSS.n1140 4.7025e+06
R19563 VSS.n1140 VSS.n1109 4.53e+06
R19564 VSS.n1106 VSS.n441 4.30038e+06
R19565 VSS.n1085 VSS.n9 3.18285e+06
R19566 VSS.n12 VSS.n11 3.11669e+06
R19567 VSS.n2913 VSS.n2912 3.1155e+06
R19568 VSS.n1135 VSS.n35 3.11369e+06
R19569 VSS.n2914 VSS.n8 3.02431e+06
R19570 VSS.n1418 VSS.n154 2.51381e+06
R19571 VSS.n2913 VSS.n10 2.499e+06
R19572 VSS.n1109 VSS.n10 2.397e+06
R19573 VSS.n1121 VSS.n11 1.68349e+06
R19574 VSS.n1135 VSS.n33 1.68349e+06
R19575 VSS.n1134 VSS.n35 1.665e+06
R19576 VSS.n2910 VSS.n12 1.662e+06
R19577 VSS.n1109 VSS.n1108 1.443e+06
R19578 VSS.n2912 VSS.n2911 1.08848e+06
R19579 VSS.n1136 VSS.n1134 1.08823e+06
R19580 VSS.n442 VSS.n441 1.044e+06
R19581 VSS.n1107 VSS.n438 1.0095e+06
R19582 VSS.n870 VSS.n416 840000
R19583 VSS.n1107 VSS.n439 815966
R19584 VSS.n1104 VSS.n442 795000
R19585 VSS.n943 VSS.n942 751088
R19586 VSS.n1136 VSS.n1135 415500
R19587 VSS.n2912 VSS.n11 415500
R19588 VSS.n1107 VSS.n1106 409562
R19589 VSS.n1107 VSS.n440 408611
R19590 VSS.n1134 VSS.n1110 277000
R19591 VSS.n2911 VSS.n7 277000
R19592 VSS.n736 VSS.n526 119767
R19593 VSS.n953 VSS.n526 102500
R19594 VSS.n582 VSS.n581 75000
R19595 VSS.n953 VSS.n491 52304.8
R19596 VSS.n1139 VSS.n1138 49582.9
R19597 VSS.n1228 VSS.n1225 48150
R19598 VSS.n872 VSS.n871 48150
R19599 VSS.n1419 VSS.n143 39237.5
R19600 VSS.n670 VSS.n601 33039.1
R19601 VSS.n841 VSS.n752 33011.2
R19602 VSS.n1254 VSS.n360 33011.2
R19603 VSS.n458 VSS.n8 31816.1
R19604 VSS.n438 VSS.n434 30464.8
R19605 VSS.n1108 VSS.n435 29621.2
R19606 VSS.n1378 VSS.n327 28106.7
R19607 VSS.n1005 VSS.n459 27000
R19608 VSS.n1005 VSS.n491 27000
R19609 VSS.n1083 VSS.n459 27000
R19610 VSS.n1111 VSS.n430 25026.3
R19611 VSS.n460 VSS.n436 24089.8
R19612 VSS.n1026 VSS.n437 24089.8
R19613 VSS.n937 VSS.n435 22834.8
R19614 VSS.n1105 VSS.n440 22334.8
R19615 VSS.n1007 VSS.n439 21736.5
R19616 VSS.n1228 VSS.n1227 21144.3
R19617 VSS.n942 VSS.n941 20874.3
R19618 VSS.n940 VSS.n491 19539
R19619 VSS.n1001 VSS.n459 19066
R19620 VSS.n941 VSS.n940 18914.1
R19621 VSS.n873 VSS.n872 18065.5
R19622 VSS.n1225 VSS.n1224 18065.5
R19623 VSS.n937 VSS.n754 16897.2
R19624 VSS.n572 VSS.n492 16670.7
R19625 VSS.n1005 VSS.n1004 15986.5
R19626 VSS.n601 VSS.n583 15936.8
R19627 VSS.n1137 VSS.n1136 15370.2
R19628 VSS.n943 VSS.n939 14914.3
R19629 VSS.n572 VSS.n8 14795.8
R19630 VSS.n582 VSS.n528 10371.7
R19631 VSS.n980 VSS.n458 9815.34
R19632 VSS.n953 VSS.n528 9144.98
R19633 VSS.n942 VSS.n438 8473.45
R19634 VSS.n1227 VSS.n154 7780.74
R19635 VSS.n669 VSS.n647 7414.81
R19636 VSS.n1093 VSS.n1085 7003.19
R19637 VSS.n1006 VSS.n1005 6755.73
R19638 VSS.n1027 VSS.n459 6755.73
R19639 VSS.n1083 VSS.n1082 6755.73
R19640 VSS.n870 VSS.n869 6749.17
R19641 VSS.n1085 VSS.n1084 6507.56
R19642 VSS.n1084 VSS.n1083 6427.48
R19643 VSS.n461 VSS.n460 6068.7
R19644 VSS.n1107 VSS.n436 6068.7
R19645 VSS.n1028 VSS.n1026 6068.7
R19646 VSS.n1008 VSS.n1007 6068.7
R19647 VSS.n1107 VSS.n437 6068.7
R19648 VSS.n492 VSS.n458 5926.03
R19649 VSS.n387 VSS.n386 5627.91
R19650 VSS.n856 VSS.n855 5627.91
R19651 VSS.n910 VSS.n909 5627.91
R19652 VSS.n1164 VSS.n1158 5627.91
R19653 VSS.n671 VSS.n607 5557.43
R19654 VSS.n1141 VSS.n430 5250
R19655 VSS.n387 VSS.n374 4711.06
R19656 VSS.n856 VSS.n819 4711.06
R19657 VSS.n909 VSS.n908 4711.06
R19658 VSS.n1162 VSS.n1158 4711.06
R19659 VSS.n388 VSS.n387 4624.2
R19660 VSS.n909 VSS.n907 4624.2
R19661 VSS.n857 VSS.n856 4624.2
R19662 VSS.n1160 VSS.n1158 4624.2
R19663 VSS.n326 VSS.n155 4526.5
R19664 VSS.n573 VSS.n572 3971.15
R19665 VSS.n1105 VSS.n1104 3958.31
R19666 VSS.n1138 VSS.n1111 3800.83
R19667 VSS.n647 VSS.n574 3575.48
R19668 VSS.n1111 VSS.n360 3353.68
R19669 VSS.n1104 VSS.n1103 3293.44
R19670 VSS.n1084 VSS.n458 2973.86
R19671 VSS.n939 VSS.n938 2851.72
R19672 VSS.n1108 VSS.n1107 2783.68
R19673 VSS.n607 VSS.n580 2681.05
R19674 VSS.n1108 VSS.n433 2648.96
R19675 VSS.n1225 VSS.n416 2172
R19676 VSS.n872 VSS.n416 2172
R19677 VSS.n939 VSS.n752 2157.5
R19678 VSS.n1001 VSS.n492 1703.92
R19679 VSS.n1140 VSS.n1139 1693.37
R19680 VSS.n1115 VSS.n10 1690.55
R19681 VSS.n1137 VSS.n1112 1670.19
R19682 VSS.n1004 VSS.n492 1277.67
R19683 VSS.n1176 VSS.n1175 1273.5
R19684 VSS.n838 VSS.n837 1271.14
R19685 VSS.n1014 VSS.n489 1155.83
R19686 VSS.n1034 VSS.n1024 1155.83
R19687 VSS.n1051 VSS.n1044 1155.83
R19688 VSS.n1079 VSS.n462 1155.83
R19689 VSS.n1139 VSS.n430 1140.49
R19690 VSS.n870 VSS.n154 1035.76
R19691 VSS.n1115 VSS.n1110 989.362
R19692 VSS.n2915 VSS.n7 835.087
R19693 VSS.n836 VSS.n754 806.716
R19694 VSS.n1157 VSS.n1156 806.716
R19695 VSS.n840 VSS.n839 806.509
R19696 VSS.n1177 VSS.n363 806.509
R19697 VSS.n1134 VSS.n1133 783.213
R19698 VSS.n2910 VSS.n2909 780.513
R19699 VSS.n847 VSS.n841 745.394
R19700 VSS.n1254 VSS.n1253 745.394
R19701 VSS.n574 VSS.n492 693.078
R19702 VSS.n1108 VSS.n434 667.145
R19703 VSS.n1103 VSS.n443 570.212
R19704 VSS.n1094 VSS.n1093 568.742
R19705 VSS.n360 VSS.n327 559.968
R19706 VSS.n752 VSS.n143 551.506
R19707 VSS.n953 VSS.n952 546.929
R19708 VSS.n2909 VSS.n13 532.101
R19709 VSS.n1133 VSS.n13 532.097
R19710 VSS.n1112 VSS.n20 483.349
R19711 VSS.n1116 VSS.n1115 483.349
R19712 VSS.n2915 VSS.n2914 468.538
R19713 VSS.n581 VSS.n580 427.767
R19714 VSS.n84 VSS.n12 414.894
R19715 VSS.n2902 VSS.n35 414.894
R19716 VSS.n2914 VSS.n2913 397.651
R19717 VSS.n2913 VSS.n9 391.414
R19718 VSS.n1221 VSS.n1220 381.036
R19719 VSS.n1233 VSS.n410 381.036
R19720 VSS.n385 VSS.n384 365.483
R19721 VSS.n376 VSS.n361 365.483
R19722 VSS.n871 VSS.n868 365.483
R19723 VSS.n850 VSS.n848 365.483
R19724 VSS.n828 VSS.n827 365.483
R19725 VSS.n916 VSS.n915 365.483
R19726 VSS.n1166 VSS.n1165 365.483
R19727 VSS.n1172 VSS.n1171 365.483
R19728 VSS.n1231 VSS.n1228 365.483
R19729 VSS.n895 VSS.n778 335.351
R19730 VSS.n798 VSS.n797 335.351
R19731 VSS.n1219 VSS.n1218 335.351
R19732 VSS.n1236 VSS.n1234 335.351
R19733 VSS.n1235 VSS.n367 319.373
R19734 VSS.n898 VSS.n776 319.373
R19735 VSS.n803 VSS.n802 319.373
R19736 VSS.n421 VSS.n420 319.373
R19737 VSS.n407 VSS.n405 312.656
R19738 VSS.n406 VSS.n369 312.656
R19739 VSS.n401 VSS.n399 312.656
R19740 VSS.n400 VSS.n371 312.656
R19741 VSS.n395 VSS.n393 312.656
R19742 VSS.n394 VSS.n390 312.656
R19743 VSS.n903 VSS.n770 312.656
R19744 VSS.n889 VSS.n886 312.656
R19745 VSS.n902 VSS.n772 312.656
R19746 VSS.n891 VSS.n884 312.656
R19747 VSS.n900 VSS.n774 312.656
R19748 VSS.n893 VSS.n882 312.656
R19749 VSS.n860 VSS.n859 312.656
R19750 VSS.n813 VSS.n790 312.656
R19751 VSS.n815 VSS.n814 312.656
R19752 VSS.n807 VSS.n792 312.656
R19753 VSS.n809 VSS.n808 312.656
R19754 VSS.n801 VSS.n794 312.656
R19755 VSS.n1210 VSS.n1208 312.656
R19756 VSS.n1209 VSS.n423 312.656
R19757 VSS.n1204 VSS.n1202 312.656
R19758 VSS.n1203 VSS.n425 312.656
R19759 VSS.n1198 VSS.n1196 312.656
R19760 VSS.n1197 VSS.n427 312.656
R19761 VSS.n583 VSS.n582 312.269
R19762 VSS.n1156 VSS.n430 306.687
R19763 VSS.n1013 VSS.n1008 281.534
R19764 VSS.n1006 VSS.n478 281.534
R19765 VSS.n1033 VSS.n1028 281.534
R19766 VSS.n1027 VSS.n470 281.534
R19767 VSS.n1050 VSS.n461 281.534
R19768 VSS.n1082 VSS.n1081 281.534
R19769 VSS.n96 VSS.n13 281.432
R19770 VSS.n28 VSS.n13 281.432
R19771 VSS.n389 VSS.n388 264.904
R19772 VSS.n1160 VSS.n1159 264.904
R19773 VSS.n855 VSS.n853 263.017
R19774 VSS.n911 VSS.n910 263.017
R19775 VSS.n907 VSS.n887 261.182
R19776 VSS.n858 VSS.n857 261.182
R19777 VSS.n848 VSS.n840 250.994
R19778 VSS.n363 VSS.n361 250.994
R19779 VSS.n386 VSS.n385 243.655
R19780 VSS.n1165 VSS.n1164 243.655
R19781 VSS.n1094 VSS.n442 236.268
R19782 VSS.n450 VSS.n442 228.189
R19783 VSS.n839 VSS.n838 219.947
R19784 VSS.n2905 VSS.n21 218.722
R19785 VSS.n31 VSS.n17 218.722
R19786 VSS.n1123 VSS.n1122 218.722
R19787 VSS.n1118 VSS.n1117 218.722
R19788 VSS.n1177 VSS.n1176 214.855
R19789 VSS.n2916 VSS.n2915 213.216
R19790 VSS.n2904 VSS.n15 207.922
R19791 VSS.n27 VSS.n19 207.922
R19792 VSS.n25 VSS.n16 207.922
R19793 VSS.n26 VSS.n18 207.922
R19794 VSS.n1125 VSS.n1124 207.922
R19795 VSS.n1129 VSS.n1128 207.922
R19796 VSS.n1127 VSS.n1126 207.922
R19797 VSS.n1120 VSS.n1119 207.922
R19798 VSS.n1162 VSS.n1161 182.382
R19799 VSS.n838 VSS.n836 173.287
R19800 VSS.n1176 VSS.n1157 168.32
R19801 VSS.n937 VSS.n936 155.988
R19802 VSS.n1140 VSS.n1110 153.942
R19803 VSS.n450 VSS.n448 152.125
R19804 VSS.n1143 VSS.n1142 134.334
R19805 VSS.n848 VSS.n847 129.114
R19806 VSS.n1253 VSS.n361 129.114
R19807 VSS.n375 VSS.n374 125.635
R19808 VSS.n854 VSS.n819 125.635
R19809 VSS.n908 VSS.n769 125.635
R19810 VSS.n1164 VSS.n1163 125.632
R19811 VSS.n374 VSS.n373 123.561
R19812 VSS.n908 VSS.n888 123.561
R19813 VSS.n819 VSS.n818 123.561
R19814 VSS.n386 VSS.n375 121.828
R19815 VSS.n737 VSS.n573 119.469
R19816 VSS.n855 VSS.n854 118.02
R19817 VSS.n910 VSS.n769 118.02
R19818 VSS.n907 VSS.n888 116.678
R19819 VSS.n857 VSS.n818 116.678
R19820 VSS.n1078 VSS.n442 113.647
R19821 VSS.n388 VSS.n373 112.957
R19822 VSS.n940 VSS.n486 112.356
R19823 VSS.n1161 VSS.n1160 107.941
R19824 VSS.n1163 VSS.n1162 93.7189
R19825 VSS.n1112 VSS.n7 93.3051
R19826 VSS.n581 VSS.n492 91.933
R19827 VSS.n954 VSS.n737 80.0919
R19828 VSS.n877 VSS.n778 77.4853
R19829 VSS.n797 VSS.n796 77.4853
R19830 VSS.n1220 VSS.n1219 76.793
R19831 VSS.n1234 VSS.n1233 76.793
R19832 VSS.n954 VSS.n953 68.5547
R19833 VSS.n390 VSS.n389 60.189
R19834 VSS.n903 VSS.n887 60.189
R19835 VSS.n860 VSS.n858 60.189
R19836 VSS.n1159 VSS.n427 60.189
R19837 VSS.n936 VSS.n935 48.1999
R19838 VSS.n2905 VSS.n2904 45.9051
R19839 VSS.n27 VSS.n15 45.9051
R19840 VSS.n25 VSS.n19 45.9051
R19841 VSS.n26 VSS.n16 45.9051
R19842 VSS.n31 VSS.n18 45.9051
R19843 VSS.n1124 VSS.n1123 45.9051
R19844 VSS.n1129 VSS.n1125 45.9051
R19845 VSS.n1128 VSS.n1127 45.9051
R19846 VSS.n1126 VSS.n1120 45.9051
R19847 VSS.n1119 VSS.n1118 45.9051
R19848 VSS.n895 VSS.n776 45.6858
R19849 VSS.n802 VSS.n798 45.6858
R19850 VSS.n1218 VSS.n420 45.6858
R19851 VSS.n1236 VSS.n1235 45.6858
R19852 VSS.n405 VSS.n367 44.6655
R19853 VSS.n407 VSS.n406 44.6655
R19854 VSS.n399 VSS.n369 44.6655
R19855 VSS.n401 VSS.n400 44.6655
R19856 VSS.n393 VSS.n371 44.6655
R19857 VSS.n395 VSS.n394 44.6655
R19858 VSS.n889 VSS.n770 44.6655
R19859 VSS.n902 VSS.n886 44.6655
R19860 VSS.n891 VSS.n772 44.6655
R19861 VSS.n900 VSS.n884 44.6655
R19862 VSS.n893 VSS.n774 44.6655
R19863 VSS.n898 VSS.n882 44.6655
R19864 VSS.n859 VSS.n790 44.6655
R19865 VSS.n815 VSS.n813 44.6655
R19866 VSS.n814 VSS.n792 44.6655
R19867 VSS.n809 VSS.n807 44.6655
R19868 VSS.n808 VSS.n794 44.6655
R19869 VSS.n803 VSS.n801 44.6655
R19870 VSS.n1208 VSS.n421 44.6655
R19871 VSS.n1210 VSS.n1209 44.6655
R19872 VSS.n1202 VSS.n423 44.6655
R19873 VSS.n1204 VSS.n1203 44.6655
R19874 VSS.n1196 VSS.n425 44.6655
R19875 VSS.n1198 VSS.n1197 44.6655
R19876 VSS.n941 VSS.n439 40.634
R19877 VSS.n938 VSS.n937 36.3099
R19878 VSS.n21 VSS.n20 35.104
R19879 VSS.n33 VSS.n17 35.104
R19880 VSS.n1122 VSS.n1121 35.104
R19881 VSS.n1117 VSS.n1116 35.104
R19882 VSS.n1106 VSS.n1105 34.3516
R19883 VSS.n326 VSS.n143 32.8363
R19884 VSS.n877 VSS.n876 31.799
R19885 VSS.n796 VSS.n784 31.799
R19886 VSS.n383 VSS.n382 31.1078
R19887 VSS.n381 VSS.n380 31.1078
R19888 VSS.n379 VSS.n378 31.1078
R19889 VSS.n876 VSS.n780 31.1078
R19890 VSS.n784 VSS.n783 31.1078
R19891 VSS.n849 VSS.n821 31.1078
R19892 VSS.n824 VSS.n823 31.1078
R19893 VSS.n852 VSS.n820 31.1078
R19894 VSS.n853 VSS.n852 31.1078
R19895 VSS.n823 VSS.n821 31.1078
R19896 VSS.n765 VSS.n764 31.1078
R19897 VSS.n767 VSS.n766 31.1078
R19898 VSS.n914 VSS.n768 31.1078
R19899 VSS.n768 VSS.n767 31.1078
R19900 VSS.n766 VSS.n765 31.1078
R19901 VSS.n1168 VSS.n1167 31.1078
R19902 VSS.n1170 VSS.n1169 31.1078
R19903 VSS.n1174 VSS.n1173 31.1078
R19904 VSS.n1169 VSS.n1168 31.1078
R19905 VSS.n1223 VSS.n1222 31.1078
R19906 VSS.n1230 VSS.n411 31.1078
R19907 VSS.n378 VSS.n377 31.1078
R19908 VSS.n380 VSS.n379 31.1078
R19909 VSS.n382 VSS.n381 31.1078
R19910 VSS.n751 VSS.n740 29.3111
R19911 VSS.n452 VSS.n443 28.6525
R19912 VSS.n453 VSS.n446 28.0068
R19913 VSS.n452 VSS.n446 28.0068
R19914 VSS.n327 VSS.n326 21.3837
R19915 VSS.n460 VSS.n440 17.9646
R19916 VSS.n1026 VSS.n436 17.9646
R19917 VSS.n1007 VSS.n437 17.9646
R19918 VSS.n1100 VSS.n449 17.0177
R19919 VSS.n1147 VSS.n432 17.001
R19920 VSS.n1152 VSS.n431 17.001
R19921 VSS.n851 VSS.n833 17.0005
R19922 VSS.n851 VSS.n828 17.0005
R19923 VSS.n851 VSS.n835 17.0005
R19924 VSS.n851 VSS.n850 17.0005
R19925 VSS.n862 VSS.n861 17.0005
R19926 VSS.n861 VSS.n798 17.0005
R19927 VSS.n861 VSS.n800 17.0005
R19928 VSS.n861 VSS.n803 17.0005
R19929 VSS.n861 VSS.n795 17.0005
R19930 VSS.n861 VSS.n794 17.0005
R19931 VSS.n861 VSS.n806 17.0005
R19932 VSS.n861 VSS.n809 17.0005
R19933 VSS.n861 VSS.n793 17.0005
R19934 VSS.n861 VSS.n792 17.0005
R19935 VSS.n861 VSS.n812 17.0005
R19936 VSS.n861 VSS.n815 17.0005
R19937 VSS.n861 VSS.n791 17.0005
R19938 VSS.n861 VSS.n790 17.0005
R19939 VSS.n861 VSS.n817 17.0005
R19940 VSS.n861 VSS.n860 17.0005
R19941 VSS.n864 VSS.n787 17.0005
R19942 VSS.n789 VSS.n788 17.0005
R19943 VSS.n802 VSS.n788 17.0005
R19944 VSS.n799 VSS.n788 17.0005
R19945 VSS.n801 VSS.n788 17.0005
R19946 VSS.n805 VSS.n788 17.0005
R19947 VSS.n808 VSS.n788 17.0005
R19948 VSS.n804 VSS.n788 17.0005
R19949 VSS.n807 VSS.n788 17.0005
R19950 VSS.n811 VSS.n788 17.0005
R19951 VSS.n814 VSS.n788 17.0005
R19952 VSS.n810 VSS.n788 17.0005
R19953 VSS.n813 VSS.n788 17.0005
R19954 VSS.n816 VSS.n788 17.0005
R19955 VSS.n859 VSS.n788 17.0005
R19956 VSS.n854 VSS.n788 17.0005
R19957 VSS.n827 VSS.n788 17.0005
R19958 VSS.n867 VSS.n785 17.0005
R19959 VSS.n868 VSS.n867 17.0005
R19960 VSS.n736 VSS.n583 17.0005
R19961 VSS.n698 VSS.n600 17.0005
R19962 VSS.n698 VSS.n601 17.0005
R19963 VSS.n673 VSS.n672 17.0005
R19964 VSS.n736 VSS.n576 17.0005
R19965 VSS.n736 VSS.n577 17.0005
R19966 VSS.n736 VSS.n578 17.0005
R19967 VSS.n736 VSS.n579 17.0005
R19968 VSS.n698 VSS.n615 17.0005
R19969 VSS.n698 VSS.n614 17.0005
R19970 VSS.n699 VSS.n698 17.0005
R19971 VSS.n698 VSS.n594 17.0005
R19972 VSS.n698 VSS.n613 17.0005
R19973 VSS.n698 VSS.n611 17.0005
R19974 VSS.n698 VSS.n609 17.0005
R19975 VSS.n698 VSS.n608 17.0005
R19976 VSS.n1002 VSS.n503 17.0005
R19977 VSS.n1002 VSS.n502 17.0005
R19978 VSS.n1002 VSS.n501 17.0005
R19979 VSS.n964 VSS.n495 17.0005
R19980 VSS.n515 VSS.n495 17.0005
R19981 VSS.n960 VSS.n959 17.0005
R19982 VSS.n959 VSS.n958 17.0005
R19983 VSS.n956 VSS.n955 17.0005
R19984 VSS.n955 VSS.n522 17.0005
R19985 VSS.n955 VSS.n528 17.0005
R19986 VSS.n955 VSS.n527 17.0005
R19987 VSS.n955 VSS.n526 17.0005
R19988 VSS.n1002 VSS.n498 17.0005
R19989 VSS.n1002 VSS.n499 17.0005
R19990 VSS.n1002 VSS.n497 17.0005
R19991 VSS.n1002 VSS.n500 17.0005
R19992 VSS.n1002 VSS.n496 17.0005
R19993 VSS.n1002 VSS.n1000 17.0005
R19994 VSS.n698 VSS.n604 17.0005
R19995 VSS.n698 VSS.n605 17.0005
R19996 VSS.n698 VSS.n603 17.0005
R19997 VSS.n698 VSS.n606 17.0005
R19998 VSS.n698 VSS.n602 17.0005
R19999 VSS.n698 VSS.n646 17.0005
R20000 VSS.n904 VSS.n896 17.0005
R20001 VSS.n904 VSS.n895 17.0005
R20002 VSS.n904 VSS.n897 17.0005
R20003 VSS.n904 VSS.n898 17.0005
R20004 VSS.n904 VSS.n894 17.0005
R20005 VSS.n904 VSS.n893 17.0005
R20006 VSS.n904 VSS.n899 17.0005
R20007 VSS.n904 VSS.n900 17.0005
R20008 VSS.n904 VSS.n892 17.0005
R20009 VSS.n904 VSS.n891 17.0005
R20010 VSS.n904 VSS.n901 17.0005
R20011 VSS.n904 VSS.n902 17.0005
R20012 VSS.n904 VSS.n890 17.0005
R20013 VSS.n904 VSS.n889 17.0005
R20014 VSS.n905 VSS.n904 17.0005
R20015 VSS.n904 VSS.n903 17.0005
R20016 VSS.n879 VSS.n878 17.0005
R20017 VSS.n921 VSS.n777 17.0005
R20018 VSS.n921 VSS.n776 17.0005
R20019 VSS.n921 VSS.n881 17.0005
R20020 VSS.n921 VSS.n882 17.0005
R20021 VSS.n921 VSS.n775 17.0005
R20022 VSS.n921 VSS.n774 17.0005
R20023 VSS.n921 VSS.n883 17.0005
R20024 VSS.n921 VSS.n884 17.0005
R20025 VSS.n921 VSS.n773 17.0005
R20026 VSS.n921 VSS.n772 17.0005
R20027 VSS.n921 VSS.n885 17.0005
R20028 VSS.n921 VSS.n886 17.0005
R20029 VSS.n921 VSS.n771 17.0005
R20030 VSS.n921 VSS.n770 17.0005
R20031 VSS.n875 VSS.n782 17.0005
R20032 VSS.n875 VSS.n873 17.0005
R20033 VSS.n912 VSS.n762 17.0005
R20034 VSS.n915 VSS.n762 17.0005
R20035 VSS.n923 VSS.n762 17.0005
R20036 VSS.n837 VSS.n762 17.0005
R20037 VSS.n921 VSS.n769 17.0005
R20038 VSS.n921 VSS.n916 17.0005
R20039 VSS.n846 VSS.n845 17.0005
R20040 VSS.n847 VSS.n846 17.0005
R20041 VSS.n929 VSS.n753 17.0005
R20042 VSS.n932 VSS.n755 17.0005
R20043 VSS.n935 VSS.n934 17.0005
R20044 VSS.n955 VSS.n529 17.0005
R20045 VSS.n955 VSS.n525 17.0005
R20046 VSS.n955 VSS.n530 17.0005
R20047 VSS.n955 VSS.n524 17.0005
R20048 VSS.n955 VSS.n571 17.0005
R20049 VSS.n698 VSS.n599 17.0005
R20050 VSS.n698 VSS.n648 17.0005
R20051 VSS.n698 VSS.n598 17.0005
R20052 VSS.n698 VSS.n649 17.0005
R20053 VSS.n698 VSS.n597 17.0005
R20054 VSS.n698 VSS.n697 17.0005
R20055 VSS.n1021 VSS.n482 17.0005
R20056 VSS.n1041 VSS.n474 17.0005
R20057 VSS.n1058 VSS.n466 17.0005
R20058 VSS.n1077 VSS.n1076 17.0005
R20059 VSS.n2903 VSS.n21 17.0005
R20060 VSS.n2903 VSS.n33 17.0005
R20061 VSS.n2903 VSS.n31 17.0005
R20062 VSS.n2903 VSS.n26 17.0005
R20063 VSS.n2903 VSS.n25 17.0005
R20064 VSS.n2903 VSS.n27 17.0005
R20065 VSS.n2904 VSS.n2903 17.0005
R20066 VSS.n2918 VSS.n2916 17.0005
R20067 VSS.n2903 VSS.n28 17.0005
R20068 VSS.n2903 VSS.n24 17.0005
R20069 VSS.n2903 VSS.n29 17.0005
R20070 VSS.n2903 VSS.n23 17.0005
R20071 VSS.n2903 VSS.n30 17.0005
R20072 VSS.n2903 VSS.n22 17.0005
R20073 VSS.n2903 VSS.n2902 17.0005
R20074 VSS.n98 VSS.n84 17.0005
R20075 VSS.n1129 VSS.n1113 17.0005
R20076 VSS.n1120 VSS.n1113 17.0005
R20077 VSS.n1118 VSS.n1113 17.0005
R20078 VSS.n1130 VSS.n1118 17.0005
R20079 VSS.n1130 VSS.n1120 17.0005
R20080 VSS.n1130 VSS.n1129 17.0005
R20081 VSS.n1121 VSS.n98 17.0005
R20082 VSS.n1123 VSS.n98 17.0005
R20083 VSS.n1125 VSS.n98 17.0005
R20084 VSS.n1128 VSS.n98 17.0005
R20085 VSS.n1126 VSS.n98 17.0005
R20086 VSS.n1119 VSS.n98 17.0005
R20087 VSS.n1117 VSS.n98 17.0005
R20088 VSS.n1181 VSS.n428 17.0005
R20089 VSS.n1172 VSS.n428 17.0005
R20090 VSS.n1189 VSS.n428 17.0005
R20091 VSS.n1166 VSS.n428 17.0005
R20092 VSS.n1175 VSS.n419 17.0005
R20093 VSS.n1171 VSS.n419 17.0005
R20094 VSS.n1165 VSS.n419 17.0005
R20095 VSS.n1217 VSS.n1192 17.0005
R20096 VSS.n1217 VSS.n427 17.0005
R20097 VSS.n1217 VSS.n1195 17.0005
R20098 VSS.n1217 VSS.n1198 17.0005
R20099 VSS.n1217 VSS.n426 17.0005
R20100 VSS.n1217 VSS.n425 17.0005
R20101 VSS.n1217 VSS.n1201 17.0005
R20102 VSS.n1217 VSS.n1204 17.0005
R20103 VSS.n1217 VSS.n424 17.0005
R20104 VSS.n1217 VSS.n423 17.0005
R20105 VSS.n1217 VSS.n1207 17.0005
R20106 VSS.n1217 VSS.n1210 17.0005
R20107 VSS.n1217 VSS.n422 17.0005
R20108 VSS.n1217 VSS.n421 17.0005
R20109 VSS.n1161 VSS.n419 17.0005
R20110 VSS.n1191 VSS.n419 17.0005
R20111 VSS.n1194 VSS.n419 17.0005
R20112 VSS.n1197 VSS.n419 17.0005
R20113 VSS.n1193 VSS.n419 17.0005
R20114 VSS.n1196 VSS.n419 17.0005
R20115 VSS.n1200 VSS.n419 17.0005
R20116 VSS.n1203 VSS.n419 17.0005
R20117 VSS.n1199 VSS.n419 17.0005
R20118 VSS.n1202 VSS.n419 17.0005
R20119 VSS.n1206 VSS.n419 17.0005
R20120 VSS.n1209 VSS.n419 17.0005
R20121 VSS.n1205 VSS.n419 17.0005
R20122 VSS.n1208 VSS.n419 17.0005
R20123 VSS.n1224 VSS.n417 17.0005
R20124 VSS.n1217 VSS.n1216 17.0005
R20125 VSS.n1218 VSS.n1217 17.0005
R20126 VSS.n1221 VSS.n418 17.0005
R20127 VSS.n1215 VSS.n419 17.0005
R20128 VSS.n420 VSS.n419 17.0005
R20129 VSS.n1214 VSS.n419 17.0005
R20130 VSS.n1213 VSS.n419 17.0005
R20131 VSS.n1232 VSS.n1231 17.0005
R20132 VSS.n1238 VSS.n1237 17.0005
R20133 VSS.n1237 VSS.n390 17.0005
R20134 VSS.n1237 VSS.n392 17.0005
R20135 VSS.n1237 VSS.n395 17.0005
R20136 VSS.n1237 VSS.n372 17.0005
R20137 VSS.n1237 VSS.n371 17.0005
R20138 VSS.n1237 VSS.n398 17.0005
R20139 VSS.n1237 VSS.n401 17.0005
R20140 VSS.n1237 VSS.n370 17.0005
R20141 VSS.n1237 VSS.n369 17.0005
R20142 VSS.n1237 VSS.n404 17.0005
R20143 VSS.n1237 VSS.n407 17.0005
R20144 VSS.n1237 VSS.n368 17.0005
R20145 VSS.n1237 VSS.n367 17.0005
R20146 VSS.n1237 VSS.n409 17.0005
R20147 VSS.n1237 VSS.n1236 17.0005
R20148 VSS.n1249 VSS.n364 17.0005
R20149 VSS.n376 VSS.n364 17.0005
R20150 VSS.n1241 VSS.n364 17.0005
R20151 VSS.n384 VSS.n364 17.0005
R20152 VSS.n1229 VSS.n410 17.0005
R20153 VSS.n385 VSS.n365 17.0005
R20154 VSS.n375 VSS.n365 17.0005
R20155 VSS.n1239 VSS.n365 17.0005
R20156 VSS.n366 VSS.n365 17.0005
R20157 VSS.n394 VSS.n365 17.0005
R20158 VSS.n391 VSS.n365 17.0005
R20159 VSS.n393 VSS.n365 17.0005
R20160 VSS.n397 VSS.n365 17.0005
R20161 VSS.n400 VSS.n365 17.0005
R20162 VSS.n396 VSS.n365 17.0005
R20163 VSS.n399 VSS.n365 17.0005
R20164 VSS.n403 VSS.n365 17.0005
R20165 VSS.n406 VSS.n365 17.0005
R20166 VSS.n402 VSS.n365 17.0005
R20167 VSS.n405 VSS.n365 17.0005
R20168 VSS.n408 VSS.n365 17.0005
R20169 VSS.n1235 VSS.n365 17.0005
R20170 VSS.n413 VSS.n365 17.0005
R20171 VSS.n414 VSS.n365 17.0005
R20172 VSS.n1252 VSS.n1251 17.0005
R20173 VSS.n1253 VSS.n1252 17.0005
R20174 VSS.n1378 VSS.n318 17.0005
R20175 VSS.n1378 VSS.n319 17.0005
R20176 VSS.n1378 VSS.n317 17.0005
R20177 VSS.n1378 VSS.n320 17.0005
R20178 VSS.n1378 VSS.n316 17.0005
R20179 VSS.n1378 VSS.n321 17.0005
R20180 VSS.n1378 VSS.n315 17.0005
R20181 VSS.n1378 VSS.n322 17.0005
R20182 VSS.n1378 VSS.n314 17.0005
R20183 VSS.n1378 VSS.n323 17.0005
R20184 VSS.n1378 VSS.n313 17.0005
R20185 VSS.n1378 VSS.n324 17.0005
R20186 VSS.n1378 VSS.n312 17.0005
R20187 VSS.n1378 VSS.n325 17.0005
R20188 VSS.n1419 VSS.n152 17.0005
R20189 VSS.n1419 VSS.n151 17.0005
R20190 VSS.n1419 VSS.n150 17.0005
R20191 VSS.n1419 VSS.n149 17.0005
R20192 VSS.n1419 VSS.n148 17.0005
R20193 VSS.n1419 VSS.n147 17.0005
R20194 VSS.n1419 VSS.n146 17.0005
R20195 VSS.n1419 VSS.n145 17.0005
R20196 VSS.n1419 VSS.n144 17.0005
R20197 VSS.n1420 VSS.n1419 17.0005
R20198 VSS.n1419 VSS.n135 17.0005
R20199 VSS.n1419 VSS.n136 17.0005
R20200 VSS.n1419 VSS.n134 17.0005
R20201 VSS.n1419 VSS.n137 17.0005
R20202 VSS.n1419 VSS.n133 17.0005
R20203 VSS.n1419 VSS.n138 17.0005
R20204 VSS.n1419 VSS.n132 17.0005
R20205 VSS.n1419 VSS.n139 17.0005
R20206 VSS.n1419 VSS.n131 17.0005
R20207 VSS.n1419 VSS.n141 17.0005
R20208 VSS.n1419 VSS.n130 17.0005
R20209 VSS.n1419 VSS.n142 17.0005
R20210 VSS.n1419 VSS.n129 17.0005
R20211 VSS.n1419 VSS.n153 17.0005
R20212 VSS.n1417 VSS.n157 17.0005
R20213 VSS.n1417 VSS.n156 17.0005
R20214 VSS.n1417 VSS.n1416 17.0005
R20215 VSS.n1386 VSS.n1385 17.0005
R20216 VSS.n1387 VSS.n1386 17.0005
R20217 VSS.n1386 VSS.n296 17.0005
R20218 VSS.n1378 VSS.n311 17.0005
R20219 VSS.n1378 VSS.n328 17.0005
R20220 VSS.n1378 VSS.n310 17.0005
R20221 VSS.n1378 VSS.n330 17.0005
R20222 VSS.n1378 VSS.n309 17.0005
R20223 VSS.n1378 VSS.n331 17.0005
R20224 VSS.n1378 VSS.n308 17.0005
R20225 VSS.n1378 VSS.n1377 17.0005
R20226 VSS.n1379 VSS.n1378 17.0005
R20227 VSS.n1378 VSS.n306 17.0005
R20228 VSS.n1145 VSS.n432 17.0005
R20229 VSS.n1150 VSS.n431 17.0005
R20230 VSS.n1100 VSS.n448 17.0005
R20231 VSS.n1097 VSS.n454 17.0005
R20232 VSS.n377 VSS.n376 15.5541
R20233 VSS.n827 VSS.n824 15.5541
R20234 VSS.n868 VSS.n783 15.5541
R20235 VSS.n828 VSS.n820 15.5541
R20236 VSS.n850 VSS.n849 15.5541
R20237 VSS.n873 VSS.n780 15.5541
R20238 VSS.n916 VSS.n914 15.5541
R20239 VSS.n915 VSS.n911 15.5541
R20240 VSS.n837 VSS.n764 15.5541
R20241 VSS.n1175 VSS.n1174 15.5541
R20242 VSS.n1171 VSS.n1170 15.5541
R20243 VSS.n1173 VSS.n1172 15.5541
R20244 VSS.n1167 VSS.n1166 15.5541
R20245 VSS.n1222 VSS.n1221 15.5541
R20246 VSS.n1224 VSS.n1223 15.5541
R20247 VSS.n411 VSS.n410 15.5541
R20248 VSS.n1231 VSS.n1230 15.5541
R20249 VSS.n384 VSS.n383 15.5541
R20250 VSS.n935 VSS.n434 15.3991
R20251 VSS.n686 VSS 14.2787
R20252 VSS.n453 VSS.n448 14.0036
R20253 VSS.n97 VSS.n96 13.72
R20254 VSS.n97 VSS.n87 13.72
R20255 VSS.n88 VSS.n85 13.6083
R20256 VSS.n90 VSS.n86 13.6083
R20257 VSS.n92 VSS.n86 13.6083
R20258 VSS.n94 VSS.n85 13.6083
R20259 VSS.n2805 VSS.n2804 12.7678
R20260 VSS.n1163 VSS.n419 12.6823
R20261 VSS.n373 VSS.n365 11.5182
R20262 VSS.n818 VSS.n788 11.5182
R20263 VSS.n921 VSS.n888 11.5182
R20264 VSS.n945 VSS.n943 11.1463
R20265 VSS.n740 VSS.n738 9.90712
R20266 VSS.n946 VSS.n751 9.24873
R20267 VSS.n656 VSS.n596 9.11426
R20268 VSS.n539 VSS.n523 9.10364
R20269 VSS.n985 VSS.n981 9.10243
R20270 VSS.n541 VSS.n539 9.08348
R20271 VSS.n1102 VSS.n1101 9.08291
R20272 VSS.n1071 VSS.n1061 9.08291
R20273 VSS.n1068 VSS.n1065 9.08291
R20274 VSS.n1053 VSS.n468 9.08291
R20275 VSS.n1048 VSS.n1047 9.08291
R20276 VSS.n1036 VSS.n476 9.08291
R20277 VSS.n1031 VSS.n1030 9.08291
R20278 VSS.n1016 VSS.n484 9.08291
R20279 VSS.n1011 VSS.n1010 9.08291
R20280 VSS.n1092 VSS.n457 9.07736
R20281 VSS.n1398 VSS.n290 9.05608
R20282 VSS.n1439 VSS.n1438 9.05608
R20283 VSS.n1312 VSS.n1311 9.05577
R20284 VSS.n2917 VSS.n4 9.04875
R20285 VSS.n746 VSS.n744 9.02498
R20286 VSS.n2876 VSS.n2875 9.02192
R20287 VSS.n635 VSS.n604 9.00165
R20288 VSS.n989 VSS.n498 9.00154
R20289 VSS.n445 VSS.n444 9.0005
R20290 VSS.n1087 VSS.n1086 9.0005
R20291 VSS.n1089 VSS.n1088 9.0005
R20292 VSS.n1091 VSS.n1090 9.0005
R20293 VSS.n1070 VSS.n1069 9.0005
R20294 VSS.n1073 VSS.n1072 9.0005
R20295 VSS.n1046 VSS.n467 9.0005
R20296 VSS.n1055 VSS.n1054 9.0005
R20297 VSS.n1029 VSS.n475 9.0005
R20298 VSS.n1038 VSS.n1037 9.0005
R20299 VSS.n1009 VSS.n483 9.0005
R20300 VSS.n1018 VSS.n1017 9.0005
R20301 VSS.n989 VSS.n988 9.0005
R20302 VSS.n991 VSS.n510 9.0005
R20303 VSS.n993 VSS.n509 9.0005
R20304 VSS.n995 VSS.n508 9.0005
R20305 VSS.n997 VSS.n507 9.0005
R20306 VSS.n998 VSS.n506 9.0005
R20307 VSS.n972 VSS.n505 9.0005
R20308 VSS.n971 VSS.n970 9.0005
R20309 VSS.n968 VSS.n512 9.0005
R20310 VSS.n966 VSS.n514 9.0005
R20311 VSS.n560 VSS.n558 9.0005
R20312 VSS.n562 VSS.n537 9.0005
R20313 VSS.n564 VSS.n536 9.0005
R20314 VSS.n566 VSS.n535 9.0005
R20315 VSS.n568 VSS.n534 9.0005
R20316 VSS.n569 VSS.n533 9.0005
R20317 VSS.n540 VSS.n532 9.0005
R20318 VSS.n702 VSS.n701 9.0005
R20319 VSS.n593 VSS.n592 9.0005
R20320 VSS.n625 VSS.n624 9.0005
R20321 VSS.n626 VSS.n617 9.0005
R20322 VSS.n644 VSS.n618 9.0005
R20323 VSS.n643 VSS.n619 9.0005
R20324 VSS.n641 VSS.n620 9.0005
R20325 VSS.n639 VSS.n621 9.0005
R20326 VSS.n637 VSS.n633 9.0005
R20327 VSS.n635 VSS.n634 9.0005
R20328 VSS.n701 VSS.n700 9.0005
R20329 VSS.n595 VSS.n593 9.0005
R20330 VSS.n624 VSS.n623 9.0005
R20331 VSS.n617 VSS.n616 9.0005
R20332 VSS.n645 VSS.n644 9.0005
R20333 VSS.n643 VSS.n642 9.0005
R20334 VSS.n641 VSS.n640 9.0005
R20335 VSS.n639 VSS.n638 9.0005
R20336 VSS.n637 VSS.n636 9.0005
R20337 VSS.n651 VSS.n650 9.0005
R20338 VSS.n696 VSS.n695 9.0005
R20339 VSS.n653 VSS.n652 9.0005
R20340 VSS.n662 VSS.n661 9.0005
R20341 VSS.n664 VSS.n663 9.0005
R20342 VSS.n666 VSS.n665 9.0005
R20343 VSS.n677 VSS.n676 9.0005
R20344 VSS.n654 VSS.n651 9.0005
R20345 VSS.n695 VSS.n694 9.0005
R20346 VSS.n655 VSS.n653 9.0005
R20347 VSS.n690 VSS.n662 9.0005
R20348 VSS.n689 VSS.n664 9.0005
R20349 VSS.n688 VSS.n666 9.0005
R20350 VSS.n677 VSS.n667 9.0005
R20351 VSS.n657 VSS.n656 9.0005
R20352 VSS.n679 VSS.n678 9.0005
R20353 VSS.n681 VSS.n680 9.0005
R20354 VSS.n610 VSS.n585 9.0005
R20355 VSS.n707 VSS.n586 9.0005
R20356 VSS.n612 VSS.n587 9.0005
R20357 VSS.n683 VSS.n679 9.0005
R20358 VSS.n682 VSS.n681 9.0005
R20359 VSS.n588 VSS.n585 9.0005
R20360 VSS.n707 VSS.n706 9.0005
R20361 VSS.n589 VSS.n587 9.0005
R20362 VSS.n733 VSS.n732 9.0005
R20363 VSS.n727 VSS.n714 9.0005
R20364 VSS.n726 VSS.n725 9.0005
R20365 VSS.n720 VSS.n717 9.0005
R20366 VSS.n724 VSS.n723 9.0005
R20367 VSS.n716 VSS.n516 9.0005
R20368 VSS.n730 VSS.n715 9.0005
R20369 VSS.n729 VSS.n728 9.0005
R20370 VSS.n719 VSS.n718 9.0005
R20371 VSS.n722 VSS.n721 9.0005
R20372 VSS.n962 VSS.n521 9.0005
R20373 VSS.n713 VSS.n584 9.0005
R20374 VSS.n713 VSS.n710 9.0005
R20375 VSS.n713 VSS.n711 9.0005
R20376 VSS.n713 VSS.n709 9.0005
R20377 VSS.n713 VSS.n712 9.0005
R20378 VSS.n532 VSS.n531 9.0005
R20379 VSS.n570 VSS.n569 9.0005
R20380 VSS.n568 VSS.n567 9.0005
R20381 VSS.n566 VSS.n565 9.0005
R20382 VSS.n564 VSS.n563 9.0005
R20383 VSS.n562 VSS.n561 9.0005
R20384 VSS.n560 VSS.n559 9.0005
R20385 VSS.n962 VSS.n957 9.0005
R20386 VSS.n962 VSS.n518 9.0005
R20387 VSS.n962 VSS.n961 9.0005
R20388 VSS.n962 VSS.n517 9.0005
R20389 VSS.n963 VSS.n962 9.0005
R20390 VSS.n966 VSS.n965 9.0005
R20391 VSS.n968 VSS.n967 9.0005
R20392 VSS.n970 VSS.n969 9.0005
R20393 VSS.n505 VSS.n504 9.0005
R20394 VSS.n999 VSS.n998 9.0005
R20395 VSS.n997 VSS.n996 9.0005
R20396 VSS.n995 VSS.n994 9.0005
R20397 VSS.n993 VSS.n992 9.0005
R20398 VSS.n991 VSS.n990 9.0005
R20399 VSS.n1309 VSS.n1304 9.0005
R20400 VSS.n1308 VSS.n1303 9.0005
R20401 VSS.n1307 VSS.n1302 9.0005
R20402 VSS.n1261 VSS.n1260 9.0005
R20403 VSS.n1322 VSS.n1321 9.0005
R20404 VSS.n1323 VSS.n1259 9.0005
R20405 VSS.n1325 VSS.n1324 9.0005
R20406 VSS.n1326 VSS.n1258 9.0005
R20407 VSS.n1328 VSS.n1327 9.0005
R20408 VSS.n1395 VSS.n292 9.0005
R20409 VSS.n1397 VSS.n1396 9.0005
R20410 VSS.n1395 VSS.n291 9.0005
R20411 VSS.n1394 VSS.n293 9.0005
R20412 VSS.n1266 VSS.n294 9.0005
R20413 VSS.n1390 VSS.n297 9.0005
R20414 VSS.n1389 VSS.n298 9.0005
R20415 VSS.n1270 VSS.n299 9.0005
R20416 VSS.n1383 VSS.n302 9.0005
R20417 VSS.n1382 VSS.n303 9.0005
R20418 VSS.n1381 VSS.n304 9.0005
R20419 VSS.n1275 VSS.n305 9.0005
R20420 VSS.n1375 VSS.n332 9.0005
R20421 VSS.n1374 VSS.n333 9.0005
R20422 VSS.n1372 VSS.n334 9.0005
R20423 VSS.n1370 VSS.n335 9.0005
R20424 VSS.n1368 VSS.n336 9.0005
R20425 VSS.n1366 VSS.n337 9.0005
R20426 VSS.n1364 VSS.n338 9.0005
R20427 VSS.n1362 VSS.n339 9.0005
R20428 VSS.n1360 VSS.n340 9.0005
R20429 VSS.n1358 VSS.n341 9.0005
R20430 VSS.n1356 VSS.n342 9.0005
R20431 VSS.n1354 VSS.n343 9.0005
R20432 VSS.n1352 VSS.n344 9.0005
R20433 VSS.n1350 VSS.n345 9.0005
R20434 VSS.n1348 VSS.n346 9.0005
R20435 VSS.n1346 VSS.n347 9.0005
R20436 VSS.n1344 VSS.n348 9.0005
R20437 VSS.n1342 VSS.n349 9.0005
R20438 VSS.n1340 VSS.n350 9.0005
R20439 VSS.n1338 VSS.n351 9.0005
R20440 VSS.n1336 VSS.n352 9.0005
R20441 VSS.n1334 VSS.n353 9.0005
R20442 VSS.n1332 VSS.n354 9.0005
R20443 VSS.n1262 VSS.n1259 9.0005
R20444 VSS.n1321 VSS.n1320 9.0005
R20445 VSS.n1263 VSS.n1261 9.0005
R20446 VSS.n1316 VSS.n1302 9.0005
R20447 VSS.n1315 VSS.n1303 9.0005
R20448 VSS.n1314 VSS.n1304 9.0005
R20449 VSS.n1306 VSS.n1305 9.0005
R20450 VSS.n1300 VSS.n1262 9.0005
R20451 VSS.n1320 VSS.n1319 9.0005
R20452 VSS.n1318 VSS.n1263 9.0005
R20453 VSS.n1317 VSS.n1316 9.0005
R20454 VSS.n1315 VSS.n1301 9.0005
R20455 VSS.n1314 VSS.n1313 9.0005
R20456 VSS.n1397 VSS.n289 9.0005
R20457 VSS.n1264 VSS.n291 9.0005
R20458 VSS.n1265 VSS.n293 9.0005
R20459 VSS.n1267 VSS.n1266 9.0005
R20460 VSS.n1268 VSS.n297 9.0005
R20461 VSS.n1269 VSS.n298 9.0005
R20462 VSS.n1271 VSS.n1270 9.0005
R20463 VSS.n1272 VSS.n302 9.0005
R20464 VSS.n1273 VSS.n303 9.0005
R20465 VSS.n1274 VSS.n304 9.0005
R20466 VSS.n1276 VSS.n1275 9.0005
R20467 VSS.n1277 VSS.n332 9.0005
R20468 VSS.n1278 VSS.n333 9.0005
R20469 VSS.n1279 VSS.n334 9.0005
R20470 VSS.n1280 VSS.n335 9.0005
R20471 VSS.n1281 VSS.n336 9.0005
R20472 VSS.n1282 VSS.n337 9.0005
R20473 VSS.n1283 VSS.n338 9.0005
R20474 VSS.n1284 VSS.n339 9.0005
R20475 VSS.n1285 VSS.n340 9.0005
R20476 VSS.n1286 VSS.n341 9.0005
R20477 VSS.n1287 VSS.n342 9.0005
R20478 VSS.n1288 VSS.n343 9.0005
R20479 VSS.n1289 VSS.n344 9.0005
R20480 VSS.n1290 VSS.n345 9.0005
R20481 VSS.n1291 VSS.n346 9.0005
R20482 VSS.n1292 VSS.n347 9.0005
R20483 VSS.n1293 VSS.n348 9.0005
R20484 VSS.n1294 VSS.n349 9.0005
R20485 VSS.n1295 VSS.n350 9.0005
R20486 VSS.n1296 VSS.n351 9.0005
R20487 VSS.n1297 VSS.n352 9.0005
R20488 VSS.n1298 VSS.n353 9.0005
R20489 VSS.n1299 VSS.n354 9.0005
R20490 VSS.n1399 VSS.n1398 9.0005
R20491 VSS.n110 VSS.n109 9.0005
R20492 VSS.n198 VSS.n113 9.0005
R20493 VSS.n199 VSS.n114 9.0005
R20494 VSS.n200 VSS.n115 9.0005
R20495 VSS.n202 VSS.n201 9.0005
R20496 VSS.n203 VSS.n118 9.0005
R20497 VSS.n204 VSS.n119 9.0005
R20498 VSS.n205 VSS.n120 9.0005
R20499 VSS.n207 VSS.n206 9.0005
R20500 VSS.n208 VSS.n123 9.0005
R20501 VSS.n209 VSS.n124 9.0005
R20502 VSS.n210 VSS.n125 9.0005
R20503 VSS.n212 VSS.n211 9.0005
R20504 VSS.n213 VSS.n197 9.0005
R20505 VSS.n215 VSS.n214 9.0005
R20506 VSS.n194 VSS.n193 9.0005
R20507 VSS.n223 VSS.n222 9.0005
R20508 VSS.n224 VSS.n192 9.0005
R20509 VSS.n226 VSS.n225 9.0005
R20510 VSS.n189 VSS.n188 9.0005
R20511 VSS.n234 VSS.n233 9.0005
R20512 VSS.n235 VSS.n187 9.0005
R20513 VSS.n237 VSS.n236 9.0005
R20514 VSS.n184 VSS.n183 9.0005
R20515 VSS.n245 VSS.n244 9.0005
R20516 VSS.n246 VSS.n182 9.0005
R20517 VSS.n248 VSS.n247 9.0005
R20518 VSS.n179 VSS.n178 9.0005
R20519 VSS.n256 VSS.n255 9.0005
R20520 VSS.n257 VSS.n177 9.0005
R20521 VSS.n259 VSS.n258 9.0005
R20522 VSS.n174 VSS.n173 9.0005
R20523 VSS.n267 VSS.n266 9.0005
R20524 VSS.n268 VSS.n172 9.0005
R20525 VSS.n271 VSS.n270 9.0005
R20526 VSS.n269 VSS.n169 9.0005
R20527 VSS.n278 VSS.n168 9.0005
R20528 VSS.n280 VSS.n279 9.0005
R20529 VSS.n281 VSS.n160 9.0005
R20530 VSS.n282 VSS.n161 9.0005
R20531 VSS.n283 VSS.n162 9.0005
R20532 VSS.n285 VSS.n284 9.0005
R20533 VSS.n286 VSS.n165 9.0005
R20534 VSS.n1405 VSS.n287 9.0005
R20535 VSS.n1404 VSS.n288 9.0005
R20536 VSS.n1403 VSS.n1400 9.0005
R20537 VSS.n1440 VSS.n1439 9.0005
R20538 VSS.n1406 VSS.n166 9.0005
R20539 VSS.n111 VSS.n110 9.0005
R20540 VSS.n1436 VSS.n113 9.0005
R20541 VSS.n1435 VSS.n114 9.0005
R20542 VSS.n1434 VSS.n115 9.0005
R20543 VSS.n201 VSS.n116 9.0005
R20544 VSS.n1430 VSS.n118 9.0005
R20545 VSS.n1429 VSS.n119 9.0005
R20546 VSS.n1428 VSS.n120 9.0005
R20547 VSS.n206 VSS.n121 9.0005
R20548 VSS.n1424 VSS.n123 9.0005
R20549 VSS.n1423 VSS.n124 9.0005
R20550 VSS.n1422 VSS.n125 9.0005
R20551 VSS.n211 VSS.n126 9.0005
R20552 VSS.n197 VSS.n196 9.0005
R20553 VSS.n217 VSS.n215 9.0005
R20554 VSS.n219 VSS.n194 9.0005
R20555 VSS.n222 VSS.n221 9.0005
R20556 VSS.n192 VSS.n191 9.0005
R20557 VSS.n228 VSS.n226 9.0005
R20558 VSS.n230 VSS.n189 9.0005
R20559 VSS.n233 VSS.n232 9.0005
R20560 VSS.n187 VSS.n186 9.0005
R20561 VSS.n239 VSS.n237 9.0005
R20562 VSS.n241 VSS.n184 9.0005
R20563 VSS.n244 VSS.n243 9.0005
R20564 VSS.n182 VSS.n181 9.0005
R20565 VSS.n250 VSS.n248 9.0005
R20566 VSS.n252 VSS.n179 9.0005
R20567 VSS.n255 VSS.n254 9.0005
R20568 VSS.n177 VSS.n176 9.0005
R20569 VSS.n261 VSS.n259 9.0005
R20570 VSS.n263 VSS.n174 9.0005
R20571 VSS.n266 VSS.n265 9.0005
R20572 VSS.n172 VSS.n171 9.0005
R20573 VSS.n273 VSS.n271 9.0005
R20574 VSS.n275 VSS.n169 9.0005
R20575 VSS.n278 VSS.n277 9.0005
R20576 VSS.n279 VSS.n159 9.0005
R20577 VSS.n1414 VSS.n160 9.0005
R20578 VSS.n1413 VSS.n161 9.0005
R20579 VSS.n1411 VSS.n162 9.0005
R20580 VSS.n284 VSS.n163 9.0005
R20581 VSS.n1407 VSS.n165 9.0005
R20582 VSS.n1406 VSS.n1405 9.0005
R20583 VSS.n1404 VSS.n167 9.0005
R20584 VSS.n1403 VSS.n1402 9.0005
R20585 VSS.n1425 VSS.n1424 9.0005
R20586 VSS.n1426 VSS.n121 9.0005
R20587 VSS.n1428 VSS.n1427 9.0005
R20588 VSS.n1429 VSS.n117 9.0005
R20589 VSS.n1431 VSS.n1430 9.0005
R20590 VSS.n1432 VSS.n116 9.0005
R20591 VSS.n1434 VSS.n1433 9.0005
R20592 VSS.n1435 VSS.n112 9.0005
R20593 VSS.n1437 VSS.n1436 9.0005
R20594 VSS.n1408 VSS.n1407 9.0005
R20595 VSS.n1409 VSS.n163 9.0005
R20596 VSS.n1411 VSS.n1410 9.0005
R20597 VSS.n1413 VSS.n1412 9.0005
R20598 VSS.n1415 VSS.n1414 9.0005
R20599 VSS.n159 VSS.n158 9.0005
R20600 VSS.n277 VSS.n276 9.0005
R20601 VSS.n275 VSS.n274 9.0005
R20602 VSS.n273 VSS.n272 9.0005
R20603 VSS.n171 VSS.n170 9.0005
R20604 VSS.n265 VSS.n264 9.0005
R20605 VSS.n263 VSS.n262 9.0005
R20606 VSS.n261 VSS.n260 9.0005
R20607 VSS.n176 VSS.n175 9.0005
R20608 VSS.n254 VSS.n253 9.0005
R20609 VSS.n252 VSS.n251 9.0005
R20610 VSS.n250 VSS.n249 9.0005
R20611 VSS.n181 VSS.n180 9.0005
R20612 VSS.n243 VSS.n242 9.0005
R20613 VSS.n241 VSS.n240 9.0005
R20614 VSS.n239 VSS.n238 9.0005
R20615 VSS.n186 VSS.n185 9.0005
R20616 VSS.n232 VSS.n231 9.0005
R20617 VSS.n230 VSS.n229 9.0005
R20618 VSS.n228 VSS.n227 9.0005
R20619 VSS.n191 VSS.n190 9.0005
R20620 VSS.n221 VSS.n220 9.0005
R20621 VSS.n219 VSS.n218 9.0005
R20622 VSS.n217 VSS.n216 9.0005
R20623 VSS.n196 VSS.n195 9.0005
R20624 VSS.n128 VSS.n126 9.0005
R20625 VSS.n1422 VSS.n1421 9.0005
R20626 VSS.n1423 VSS.n122 9.0005
R20627 VSS.n1074 VSS.n1067 9.0005
R20628 VSS.n1056 VSS.n465 9.0005
R20629 VSS.n1039 VSS.n473 9.0005
R20630 VSS.n1019 VSS.n481 9.0005
R20631 VSS.n1021 VSS.n1020 9.0005
R20632 VSS.n1041 VSS.n1040 9.0005
R20633 VSS.n1058 VSS.n1057 9.0005
R20634 VSS.n1076 VSS.n1075 9.0005
R20635 VSS.n744 VSS.n741 9.0005
R20636 VSS.n743 VSS.n742 9.0005
R20637 VSS.n750 VSS.n749 9.0005
R20638 VSS.n745 VSS.n743 9.0005
R20639 VSS.n749 VSS.n748 9.0005
R20640 VSS.n748 VSS.n747 9.0005
R20641 VSS.n2807 VSS.n2806 9.0005
R20642 VSS.n103 VSS.n102 9.0005
R20643 VSS.n2814 VSS.n2813 9.0005
R20644 VSS.n2815 VSS.n101 9.0005
R20645 VSS.n2817 VSS.n2816 9.0005
R20646 VSS.n82 VSS.n81 9.0005
R20647 VSS.n2825 VSS.n2824 9.0005
R20648 VSS.n2826 VSS.n80 9.0005
R20649 VSS.n2828 VSS.n2827 9.0005
R20650 VSS.n76 VSS.n75 9.0005
R20651 VSS.n2836 VSS.n2835 9.0005
R20652 VSS.n2837 VSS.n74 9.0005
R20653 VSS.n2839 VSS.n2838 9.0005
R20654 VSS.n66 VSS.n65 9.0005
R20655 VSS.n2847 VSS.n2846 9.0005
R20656 VSS.n2848 VSS.n64 9.0005
R20657 VSS.n2851 VSS.n2850 9.0005
R20658 VSS.n2849 VSS.n60 9.0005
R20659 VSS.n2857 VSS.n59 9.0005
R20660 VSS.n2859 VSS.n2858 9.0005
R20661 VSS.n2860 VSS.n42 9.0005
R20662 VSS.n2861 VSS.n43 9.0005
R20663 VSS.n2862 VSS.n44 9.0005
R20664 VSS.n2864 VSS.n2863 9.0005
R20665 VSS.n2865 VSS.n48 9.0005
R20666 VSS.n2866 VSS.n49 9.0005
R20667 VSS.n2867 VSS.n50 9.0005
R20668 VSS.n2868 VSS.n51 9.0005
R20669 VSS.n2869 VSS.n52 9.0005
R20670 VSS.n2871 VSS.n2870 9.0005
R20671 VSS.n2872 VSS.n55 9.0005
R20672 VSS.n2873 VSS.n56 9.0005
R20673 VSS.n2874 VSS.n57 9.0005
R20674 VSS.n2805 VSS.n107 9.0005
R20675 VSS.n2808 VSS.n2807 9.0005
R20676 VSS.n104 VSS.n103 9.0005
R20677 VSS.n2813 VSS.n2812 9.0005
R20678 VSS.n101 VSS.n100 9.0005
R20679 VSS.n2818 VSS.n2817 9.0005
R20680 VSS.n83 VSS.n82 9.0005
R20681 VSS.n2824 VSS.n2823 9.0005
R20682 VSS.n80 VSS.n79 9.0005
R20683 VSS.n2829 VSS.n2828 9.0005
R20684 VSS.n77 VSS.n76 9.0005
R20685 VSS.n2835 VSS.n2834 9.0005
R20686 VSS.n74 VSS.n73 9.0005
R20687 VSS.n2840 VSS.n2839 9.0005
R20688 VSS.n67 VSS.n66 9.0005
R20689 VSS.n2846 VSS.n2845 9.0005
R20690 VSS.n64 VSS.n63 9.0005
R20691 VSS.n2852 VSS.n2851 9.0005
R20692 VSS.n61 VSS.n60 9.0005
R20693 VSS.n2857 VSS.n2856 9.0005
R20694 VSS.n2858 VSS.n41 9.0005
R20695 VSS.n2898 VSS.n42 9.0005
R20696 VSS.n2897 VSS.n43 9.0005
R20697 VSS.n2896 VSS.n44 9.0005
R20698 VSS.n2863 VSS.n45 9.0005
R20699 VSS.n2892 VSS.n48 9.0005
R20700 VSS.n2891 VSS.n49 9.0005
R20701 VSS.n2890 VSS.n50 9.0005
R20702 VSS.n2887 VSS.n51 9.0005
R20703 VSS.n2886 VSS.n52 9.0005
R20704 VSS.n2870 VSS.n53 9.0005
R20705 VSS.n2882 VSS.n55 9.0005
R20706 VSS.n2881 VSS.n56 9.0005
R20707 VSS.n2880 VSS.n57 9.0005
R20708 VSS.n2877 VSS.n58 9.0005
R20709 VSS.n107 VSS.n106 9.0005
R20710 VSS.n2876 VSS.n14 9.0005
R20711 VSS.n2878 VSS.n2877 9.0005
R20712 VSS.n2880 VSS.n2879 9.0005
R20713 VSS.n2881 VSS.n54 9.0005
R20714 VSS.n2883 VSS.n2882 9.0005
R20715 VSS.n2884 VSS.n53 9.0005
R20716 VSS.n2886 VSS.n2885 9.0005
R20717 VSS.n2888 VSS.n2887 9.0005
R20718 VSS.n2890 VSS.n2889 9.0005
R20719 VSS.n2891 VSS.n47 9.0005
R20720 VSS.n2893 VSS.n2892 9.0005
R20721 VSS.n2894 VSS.n45 9.0005
R20722 VSS.n2896 VSS.n2895 9.0005
R20723 VSS.n2897 VSS.n40 9.0005
R20724 VSS.n2899 VSS.n2898 9.0005
R20725 VSS.n41 VSS.n39 9.0005
R20726 VSS.n2856 VSS.n2855 9.0005
R20727 VSS.n2854 VSS.n61 9.0005
R20728 VSS.n2853 VSS.n2852 9.0005
R20729 VSS.n63 VSS.n62 9.0005
R20730 VSS.n2845 VSS.n2844 9.0005
R20731 VSS.n2842 VSS.n67 9.0005
R20732 VSS.n2841 VSS.n2840 9.0005
R20733 VSS.n2832 VSS.n73 9.0005
R20734 VSS.n2834 VSS.n2833 9.0005
R20735 VSS.n2831 VSS.n77 9.0005
R20736 VSS.n2830 VSS.n2829 9.0005
R20737 VSS.n79 VSS.n78 9.0005
R20738 VSS.n2823 VSS.n2822 9.0005
R20739 VSS.n2820 VSS.n83 9.0005
R20740 VSS.n2819 VSS.n2818 9.0005
R20741 VSS.n100 VSS.n99 9.0005
R20742 VSS.n2812 VSS.n2811 9.0005
R20743 VSS.n2810 VSS.n104 9.0005
R20744 VSS.n2809 VSS.n2808 9.0005
R20745 VSS.n106 VSS.n105 9.0005
R20746 VSS.n2924 VSS.n2923 9.0005
R20747 VSS.n6 VSS.n5 9.0005
R20748 VSS.n2923 VSS.n2922 9.0005
R20749 VSS.n2919 VSS.n6 9.0005
R20750 VSS.n2922 VSS.n2921 9.0005
R20751 VSS.n2918 VSS.n2917 9.0005
R20752 VSS.n1329 VSS.n355 9.0005
R20753 VSS.n1332 VSS.n1331 9.0005
R20754 VSS.n1334 VSS.n1333 9.0005
R20755 VSS.n1336 VSS.n1335 9.0005
R20756 VSS.n1338 VSS.n1337 9.0005
R20757 VSS.n1340 VSS.n1339 9.0005
R20758 VSS.n1342 VSS.n1341 9.0005
R20759 VSS.n1344 VSS.n1343 9.0005
R20760 VSS.n1346 VSS.n1345 9.0005
R20761 VSS.n1348 VSS.n1347 9.0005
R20762 VSS.n1350 VSS.n1349 9.0005
R20763 VSS.n1352 VSS.n1351 9.0005
R20764 VSS.n1354 VSS.n1353 9.0005
R20765 VSS.n1356 VSS.n1355 9.0005
R20766 VSS.n1358 VSS.n1357 9.0005
R20767 VSS.n1360 VSS.n1359 9.0005
R20768 VSS.n1362 VSS.n1361 9.0005
R20769 VSS.n1364 VSS.n1363 9.0005
R20770 VSS.n1366 VSS.n1365 9.0005
R20771 VSS.n1368 VSS.n1367 9.0005
R20772 VSS.n1370 VSS.n1369 9.0005
R20773 VSS.n1372 VSS.n1371 9.0005
R20774 VSS.n1374 VSS.n1373 9.0005
R20775 VSS.n1376 VSS.n1375 9.0005
R20776 VSS.n307 VSS.n305 9.0005
R20777 VSS.n1381 VSS.n1380 9.0005
R20778 VSS.n1382 VSS.n301 9.0005
R20779 VSS.n1384 VSS.n1383 9.0005
R20780 VSS.n300 VSS.n299 9.0005
R20781 VSS.n1389 VSS.n1388 9.0005
R20782 VSS.n1391 VSS.n1390 9.0005
R20783 VSS.n1392 VSS.n294 9.0005
R20784 VSS.n1394 VSS.n1393 9.0005
R20785 VSS.n984 VSS.n983 9.0005
R20786 VSS.n982 VSS.n1 9.0005
R20787 VSS.n4295 VSS.n4294 9.0005
R20788 VSS.n984 VSS.n979 9.0005
R20789 VSS.n2 VSS.n1 9.0005
R20790 VSS.n4294 VSS.n4293 9.0005
R20791 VSS.n986 VSS.n985 9.0005
R20792 VSS.n542 VSS.n533 9.0005
R20793 VSS.n543 VSS.n534 9.0005
R20794 VSS.n544 VSS.n535 9.0005
R20795 VSS.n545 VSS.n536 9.0005
R20796 VSS.n546 VSS.n537 9.0005
R20797 VSS.n558 VSS.n557 9.0005
R20798 VSS.n556 VSS.n538 9.0005
R20799 VSS.n555 VSS.n554 9.0005
R20800 VSS.n553 VSS.n552 9.0005
R20801 VSS.n551 VSS.n550 9.0005
R20802 VSS.n549 VSS.n521 9.0005
R20803 VSS.n548 VSS.n514 9.0005
R20804 VSS.n547 VSS.n512 9.0005
R20805 VSS.n971 VSS.n511 9.0005
R20806 VSS.n973 VSS.n972 9.0005
R20807 VSS.n974 VSS.n506 9.0005
R20808 VSS.n975 VSS.n507 9.0005
R20809 VSS.n976 VSS.n508 9.0005
R20810 VSS.n977 VSS.n509 9.0005
R20811 VSS.n978 VSS.n510 9.0005
R20812 VSS.n988 VSS.n987 9.0005
R20813 VSS.n659 VSS.n654 9.0005
R20814 VSS.n694 VSS.n693 9.0005
R20815 VSS.n692 VSS.n655 9.0005
R20816 VSS.n691 VSS.n690 9.0005
R20817 VSS.n689 VSS.n660 9.0005
R20818 VSS.n688 VSS.n687 9.0005
R20819 VSS.n685 VSS.n667 9.0005
R20820 VSS.n684 VSS.n683 9.0005
R20821 VSS.n682 VSS.n675 9.0005
R20822 VSS.n590 VSS.n588 9.0005
R20823 VSS.n706 VSS.n705 9.0005
R20824 VSS.n704 VSS.n589 9.0005
R20825 VSS.n703 VSS.n702 9.0005
R20826 VSS.n592 VSS.n591 9.0005
R20827 VSS.n625 VSS.n622 9.0005
R20828 VSS.n627 VSS.n626 9.0005
R20829 VSS.n628 VSS.n618 9.0005
R20830 VSS.n629 VSS.n619 9.0005
R20831 VSS.n630 VSS.n620 9.0005
R20832 VSS.n631 VSS.n621 9.0005
R20833 VSS.n633 VSS.n632 9.0005
R20834 VSS.n634 VSS.n3 9.0005
R20835 VSS.n658 VSS.n657 9.0005
R20836 VSS.n1004 VSS.n494 8.501
R20837 VSS.n1004 VSS.n493 8.501
R20838 VSS.n1127 VSS.n1114 8.501
R20839 VSS.n451 VSS.n450 8.501
R20840 VSS.n757 VSS.n435 8.5005
R20841 VSS.n952 VSS.n951 8.5005
R20842 VSS.n2906 VSS.n20 8.5005
R20843 VSS.n2906 VSS.n17 8.5005
R20844 VSS.n2906 VSS.n18 8.5005
R20845 VSS.n2906 VSS.n16 8.5005
R20846 VSS.n2906 VSS.n19 8.5005
R20847 VSS.n2906 VSS.n15 8.5005
R20848 VSS.n2906 VSS.n2905 8.5005
R20849 VSS.n71 VSS.n28 8.5005
R20850 VSS.n2902 VSS.n2901 8.5005
R20851 VSS.n96 VSS.n68 8.5005
R20852 VSS.n95 VSS.n84 8.5005
R20853 VSS.n96 VSS.n95 8.5005
R20854 VSS.n95 VSS.n87 8.5005
R20855 VSS.n95 VSS.n90 8.5005
R20856 VSS.n95 VSS.n92 8.5005
R20857 VSS.n95 VSS.n88 8.5005
R20858 VSS.n95 VSS.n94 8.5005
R20859 VSS.n1122 VSS.n1113 8.5005
R20860 VSS.n1116 VSS.n1113 8.5005
R20861 VSS.n1124 VSS.n1113 8.5005
R20862 VSS.n1256 VSS.n1255 8.5005
R20863 VSS.n757 VSS.n433 8.5005
R20864 VSS.n846 VSS.n842 8.49541
R20865 VSS.n1255 VSS.n359 8.49541
R20866 VSS.n1252 VSS.n362 8.49541
R20867 VSS.n1419 VSS.n140 8.48944
R20868 VSS.n1378 VSS.n329 8.48944
R20869 VSS.n851 VSS.n830 8.48603
R20870 VSS.n851 VSS.n826 8.48603
R20871 VSS.n851 VSS.n822 8.48603
R20872 VSS.n787 VSS.n786 8.48603
R20873 VSS.n865 VSS.n787 8.48603
R20874 VSS.n863 VSS.n788 8.48603
R20875 VSS.n832 VSS.n788 8.48603
R20876 VSS.n829 VSS.n788 8.48603
R20877 VSS.n825 VSS.n788 8.48603
R20878 VSS.n834 VSS.n788 8.48603
R20879 VSS.n867 VSS.n866 8.48603
R20880 VSS.n878 VSS.n781 8.48603
R20881 VSS.n878 VSS.n779 8.48603
R20882 VSS.n921 VSS.n880 8.48603
R20883 VSS.n875 VSS.n874 8.48603
R20884 VSS.n917 VSS.n762 8.48603
R20885 VSS.n919 VSS.n762 8.48603
R20886 VSS.n763 VSS.n762 8.48603
R20887 VSS.n921 VSS.n913 8.48603
R20888 VSS.n921 VSS.n918 8.48603
R20889 VSS.n921 VSS.n920 8.48603
R20890 VSS.n922 VSS.n921 8.48603
R20891 VSS.n1183 VSS.n428 8.48603
R20892 VSS.n1185 VSS.n428 8.48603
R20893 VSS.n1187 VSS.n428 8.48603
R20894 VSS.n1182 VSS.n419 8.48603
R20895 VSS.n1184 VSS.n419 8.48603
R20896 VSS.n1186 VSS.n419 8.48603
R20897 VSS.n1188 VSS.n419 8.48603
R20898 VSS.n1212 VSS.n417 8.48603
R20899 VSS.n1232 VSS.n415 8.48603
R20900 VSS.n1247 VSS.n364 8.48603
R20901 VSS.n1245 VSS.n364 8.48603
R20902 VSS.n1243 VSS.n364 8.48603
R20903 VSS.n1248 VSS.n365 8.48603
R20904 VSS.n1246 VSS.n365 8.48603
R20905 VSS.n1244 VSS.n365 8.48603
R20906 VSS.n1242 VSS.n365 8.48603
R20907 VSS.n1095 VSS.n456 8.4728
R20908 VSS.n934 VSS.n933 8.47111
R20909 VSS.n2920 VSS.n2916 8.47111
R20910 VSS.n1077 VSS.n1066 8.4706
R20911 VSS.n466 VSS.n464 8.4706
R20912 VSS.n474 VSS.n472 8.4706
R20913 VSS.n482 VSS.n480 8.4706
R20914 VSS.n1100 VSS.n447 8.4706
R20915 VSS.n955 VSS.n523 8.44994
R20916 VSS.n698 VSS.n596 8.44466
R20917 VSS.n38 VSS.n28 7.59315
R20918 VSS.n38 VSS.n24 7.59315
R20919 VSS.n93 VSS.n84 7.55879
R20920 VSS.n91 VSS.n88 7.55879
R20921 VSS.n90 VSS.n89 7.55879
R20922 VSS.n70 VSS.n29 7.55879
R20923 VSS.n37 VSS.n23 7.55879
R20924 VSS.n69 VSS.n30 7.55879
R20925 VSS.n36 VSS.n22 7.55879
R20926 VSS.n2902 VSS.n34 7.55879
R20927 VSS.n69 VSS.n23 7.55879
R20928 VSS.n34 VSS.n22 7.55879
R20929 VSS.n70 VSS.n24 7.55879
R20930 VSS.n37 VSS.n29 7.55879
R20931 VSS.n36 VSS.n30 7.55879
R20932 VSS.n89 VSS.n87 7.55879
R20933 VSS.n92 VSS.n91 7.55879
R20934 VSS.n94 VSS.n93 7.55879
R20935 VSS.n1211 VSS.n417 5.66867
R20936 VSS.n1232 VSS.n412 5.66867
R20937 VSS.n1211 VSS.n418 5.66811
R20938 VSS.n1229 VSS.n412 5.66811
R20939 VSS.n1418 VSS.n1417 5.66717
R20940 VSS.n1386 VSS.n155 5.66717
R20941 VSS.n1255 VSS.n356 5.65785
R20942 VSS.n1095 VSS.n457 5.63627
R20943 VSS.n1080 VSS.n1062 5.63396
R20944 VSS.n1052 VSS.n469 5.63396
R20945 VSS.n1035 VSS.n477 5.63396
R20946 VSS.n1015 VSS.n485 5.63396
R20947 VSS.n1101 VSS.n1100 5.63382
R20948 VSS.n1080 VSS.n1061 5.63382
R20949 VSS.n1077 VSS.n1065 5.63382
R20950 VSS.n1053 VSS.n1052 5.63382
R20951 VSS.n1047 VSS.n466 5.63382
R20952 VSS.n1036 VSS.n1035 5.63382
R20953 VSS.n1030 VSS.n474 5.63382
R20954 VSS.n1016 VSS.n1015 5.63382
R20955 VSS.n1010 VSS.n482 5.63382
R20956 VSS.n759 VSS.n756 5.6156
R20957 VSS.n1025 VSS.n476 5.40173
R20958 VSS.n1112 VSS.n13 5.40104
R20959 VSS.n1115 VSS.n13 5.40104
R20960 VSS.n1103 VSS.n1102 5.39593
R20961 VSS.n490 VSS.n484 5.39516
R20962 VSS.n1045 VSS.n468 5.39516
R20963 VSS.n1071 VSS.n463 5.39513
R20964 VSS.n1093 VSS.n1092 5.36621
R20965 VSS.n1012 VSS.n1011 5.3654
R20966 VSS.n1032 VSS.n1031 5.3654
R20967 VSS.n1049 VSS.n1048 5.3654
R20968 VSS.n1068 VSS.n1063 5.3654
R20969 VSS.n489 VSS.n486 5.16623
R20970 VSS.n1014 VSS.n1013 5.16623
R20971 VSS.n1024 VSS.n478 5.16623
R20972 VSS.n1034 VSS.n1033 5.16623
R20973 VSS.n1044 VSS.n470 5.16623
R20974 VSS.n1051 VSS.n1050 5.16623
R20975 VSS.n1081 VSS.n462 5.16623
R20976 VSS.n1079 VSS.n1078 5.16623
R20977 VSS.n926 VSS.n754 4.76027
R20978 VSS.n1156 VSS.n1155 4.76027
R20979 VSS.n981 VSS.n980 4.69919
R20980 VSS.n292 VSS.n290 4.64528
R20981 VSS.n1310 VSS.n1309 4.64528
R20982 VSS.n1401 VSS.n166 4.64528
R20983 VSS.n1438 VSS.n1437 4.64528
R20984 VSS.n980 VSS.n0 4.58034
R20985 VSS.n542 VSS.n541 4.52011
R20986 VSS.n1313 VSS.n1312 4.5158
R20987 VSS.n747 VSS.n746 4.48901
R20988 VSS.n2924 VSS.n4 4.47713
R20989 VSS.n962 VSS.n520 4.45987
R20990 VSS.n962 VSS.n519 4.45987
R20991 VSS.n1227 VSS.n1226 4.32947
R20992 VSS.n1004 VSS.n1003 4.251
R20993 VSS.n756 VSS.n435 4.251
R20994 VSS.n758 VSS.n757 4.17719
R20995 VSS.n1008 VSS.n1006 3.8748
R20996 VSS.n1028 VSS.n1027 3.8748
R20997 VSS.n1082 VSS.n461 3.8748
R20998 VSS.n1144 VSS.n1143 3.65859
R20999 VSS.n1099 VSS.n1098 3.57718
R21000 VSS.n671 VSS.n669 3.41008
R21001 VSS.n736 VSS.n574 3.4005
R21002 VSS.n945 VSS.n944 3.1511
R21003 VSS.n947 VSS.n750 3.12829
R21004 VSS.n946 VSS.n945 3.03683
R21005 VSS.n1015 VSS.n488 2.95625
R21006 VSS.n1035 VSS.n1023 2.95625
R21007 VSS.n1052 VSS.n1043 2.95625
R21008 VSS.n1080 VSS.n1060 2.95625
R21009 VSS.n487 VSS.n482 2.9562
R21010 VSS.n479 VSS.n474 2.9562
R21011 VSS.n471 VSS.n466 2.9562
R21012 VSS.n1077 VSS.n1064 2.9562
R21013 VSS.n951 VSS.n950 2.9539
R21014 VSS.n947 VSS.n738 2.83458
R21015 VSS.n1002 VSS.n1001 2.83383
R21016 VSS.n698 VSS.n647 2.83383
R21017 VSS.n1014 VSS.n490 2.83383
R21018 VSS.n490 VSS.n486 2.83383
R21019 VSS.n1034 VSS.n1025 2.83383
R21020 VSS.n1025 VSS.n478 2.83383
R21021 VSS.n1051 VSS.n1045 2.83383
R21022 VSS.n1045 VSS.n470 2.83383
R21023 VSS.n1079 VSS.n463 2.83383
R21024 VSS.n1081 VSS.n463 2.83383
R21025 VSS.n1013 VSS.n1012 2.83383
R21026 VSS.n1012 VSS.n489 2.83383
R21027 VSS.n1033 VSS.n1032 2.83383
R21028 VSS.n1032 VSS.n1024 2.83383
R21029 VSS.n1050 VSS.n1049 2.83383
R21030 VSS.n1049 VSS.n1044 2.83383
R21031 VSS.n1078 VSS.n1063 2.83383
R21032 VSS.n1063 VSS.n462 2.83383
R21033 VSS.n1015 VSS.n486 2.83383
R21034 VSS.n1035 VSS.n478 2.83383
R21035 VSS.n1052 VSS.n470 2.83383
R21036 VSS.n1081 VSS.n1080 2.83383
R21037 VSS.n1080 VSS.n1079 2.83383
R21038 VSS.n1052 VSS.n1051 2.83383
R21039 VSS.n1035 VSS.n1034 2.83383
R21040 VSS.n1015 VSS.n1014 2.83383
R21041 VSS.n489 VSS.n482 2.83383
R21042 VSS.n1013 VSS.n482 2.83383
R21043 VSS.n1024 VSS.n474 2.83383
R21044 VSS.n1033 VSS.n474 2.83383
R21045 VSS.n1044 VSS.n466 2.83383
R21046 VSS.n1050 VSS.n466 2.83383
R21047 VSS.n1077 VSS.n462 2.83383
R21048 VSS.n1078 VSS.n1077 2.83383
R21049 VSS.n947 VSS.n946 2.83383
R21050 VSS.n948 VSS.n947 2.80958
R21051 VSS.n951 VSS.n739 2.73145
R21052 VSS.n1149 VSS.n432 2.72142
R21053 VSS.n1154 VSS.n431 2.72142
R21054 VSS.n1132 VSS.n1131 2.7174
R21055 VSS.n2911 VSS.n2910 2.70077
R21056 VSS.n944 VSS.n739 2.6007
R21057 VSS.n1096 VSS.n1095 2.48061
R21058 VSS.n955 VSS.n954 2.42907
R21059 VSS.n737 VSS.n736 2.42907
R21060 VSS.n844 VSS.n841 2.40513
R21061 VSS.n927 VSS.n753 2.30109
R21062 VSS.n930 VSS.n755 2.30109
R21063 VSS.n2939 VSS.n2925 2.2505
R21064 VSS.n4267 VSS.n4266 2.2505
R21065 VSS.n4262 VSS.n2953 2.2505
R21066 VSS.n4260 VSS.n2955 2.2505
R21067 VSS.n4256 VSS.n2958 2.2505
R21068 VSS.n4254 VSS.n2960 2.2505
R21069 VSS.n3463 VSS.n3197 2.2505
R21070 VSS.n3461 VSS.n3199 2.2505
R21071 VSS.n3457 VSS.n3202 2.2505
R21072 VSS.n3455 VSS.n3204 2.2505
R21073 VSS.n3451 VSS.n3207 2.2505
R21074 VSS.n3449 VSS.n3209 2.2505
R21075 VSS.n3384 VSS.n2926 2.2505
R21076 VSS.n3860 VSS.n3005 2.2505
R21077 VSS.n3851 VSS.n3008 2.2505
R21078 VSS.n3022 VSS.n3018 2.2505
R21079 VSS.n3826 VSS.n3020 2.2505
R21080 VSS.n3035 VSS.n3029 2.2505
R21081 VSS.n3793 VSS.n3034 2.2505
R21082 VSS.n3785 VSS.n3037 2.2505
R21083 VSS.n3782 VSS.n3781 2.2505
R21084 VSS.n3777 VSS.n3776 2.2505
R21085 VSS.n3063 VSS.n3059 2.2505
R21086 VSS.n3746 VSS.n3062 2.2505
R21087 VSS.n3734 VSS.n3065 2.2505
R21088 VSS.n3726 VSS.n3725 2.2505
R21089 VSS.n3720 VSS.n3719 2.2505
R21090 VSS.n3696 VSS.n3695 2.2505
R21091 VSS.n4198 VSS.n3005 2.2505
R21092 VSS.n3008 VSS.n3007 2.2505
R21093 VSS.n3841 VSS.n3018 2.2505
R21094 VSS.n3020 VSS.n3019 2.2505
R21095 VSS.n3806 VSS.n3035 2.2505
R21096 VSS.n3803 VSS.n3034 2.2505
R21097 VSS.n3037 VSS.n3036 2.2505
R21098 VSS.n3781 VSS.n3780 2.2505
R21099 VSS.n3778 VSS.n3777 2.2505
R21100 VSS.n3756 VSS.n3063 2.2505
R21101 VSS.n3755 VSS.n3062 2.2505
R21102 VSS.n3065 VSS.n3064 2.2505
R21103 VSS.n3725 VSS.n3724 2.2505
R21104 VSS.n3721 VSS.n3720 2.2505
R21105 VSS.n3695 VSS.n3694 2.2505
R21106 VSS.n3692 VSS.n3691 2.2505
R21107 VSS.n3091 VSS.n3090 2.2505
R21108 VSS.n3676 VSS.n3675 2.2505
R21109 VSS.n3674 VSS.n3098 2.2505
R21110 VSS.n3673 VSS.n3672 2.2505
R21111 VSS.n3100 VSS.n3099 2.2505
R21112 VSS.n3629 VSS.n3628 2.2505
R21113 VSS.n3630 VSS.n3627 2.2505
R21114 VSS.n3631 VSS.n3626 2.2505
R21115 VSS.n3625 VSS.n3115 2.2505
R21116 VSS.n3624 VSS.n3623 2.2505
R21117 VSS.n3117 VSS.n3116 2.2505
R21118 VSS.n3588 VSS.n3587 2.2505
R21119 VSS.n3595 VSS.n3586 2.2505
R21120 VSS.n3596 VSS.n3585 2.2505
R21121 VSS.n3584 VSS.n3133 2.2505
R21122 VSS.n3583 VSS.n3582 2.2505
R21123 VSS.n3135 VSS.n3134 2.2505
R21124 VSS.n3566 VSS.n3565 2.2505
R21125 VSS.n3564 VSS.n3150 2.2505
R21126 VSS.n3563 VSS.n3562 2.2505
R21127 VSS.n3152 VSS.n3151 2.2505
R21128 VSS.n3522 VSS.n3521 2.2505
R21129 VSS.n3529 VSS.n3520 2.2505
R21130 VSS.n3530 VSS.n3519 2.2505
R21131 VSS.n3518 VSS.n3169 2.2505
R21132 VSS.n3517 VSS.n3516 2.2505
R21133 VSS.n3171 VSS.n3170 2.2505
R21134 VSS.n3495 VSS.n3494 2.2505
R21135 VSS.n3493 VSS.n3182 2.2505
R21136 VSS.n3492 VSS.n3491 2.2505
R21137 VSS.n3184 VSS.n3183 2.2505
R21138 VSS.n3468 VSS.n3467 2.2505
R21139 VSS.n3469 VSS.n3466 2.2505
R21140 VSS.n3470 VSS.n3469 2.2505
R21141 VSS.n3468 VSS.n3188 2.2505
R21142 VSS.n3482 VSS.n3184 2.2505
R21143 VSS.n3491 VSS.n3490 2.2505
R21144 VSS.n3186 VSS.n3182 2.2505
R21145 VSS.n3496 VSS.n3495 2.2505
R21146 VSS.n3507 VSS.n3171 2.2505
R21147 VSS.n3516 VSS.n3515 2.2505
R21148 VSS.n3169 VSS.n3166 2.2505
R21149 VSS.n3531 VSS.n3530 2.2505
R21150 VSS.n3529 VSS.n3528 2.2505
R21151 VSS.n3522 VSS.n3157 2.2505
R21152 VSS.n3544 VSS.n3152 2.2505
R21153 VSS.n3562 VSS.n3561 2.2505
R21154 VSS.n3550 VSS.n3150 2.2505
R21155 VSS.n3567 VSS.n3566 2.2505
R21156 VSS.n3569 VSS.n3135 2.2505
R21157 VSS.n3582 VSS.n3581 2.2505
R21158 VSS.n3137 VSS.n3133 2.2505
R21159 VSS.n3597 VSS.n3596 2.2505
R21160 VSS.n3595 VSS.n3594 2.2505
R21161 VSS.n3591 VSS.n3588 2.2505
R21162 VSS.n3608 VSS.n3117 2.2505
R21163 VSS.n3623 VSS.n3622 2.2505
R21164 VSS.n3614 VSS.n3115 2.2505
R21165 VSS.n3632 VSS.n3631 2.2505
R21166 VSS.n3630 VSS.n3110 2.2505
R21167 VSS.n3629 VSS.n3107 2.2505
R21168 VSS.n3648 VSS.n3100 2.2505
R21169 VSS.n3672 VSS.n3671 2.2505
R21170 VSS.n3655 VSS.n3098 2.2505
R21171 VSS.n3677 VSS.n3676 2.2505
R21172 VSS.n3679 VSS.n3091 2.2505
R21173 VSS.n3691 VSS.n3690 2.2505
R21174 VSS.n4250 VSS.n2963 2.2505
R21175 VSS.n4249 VSS.n2964 2.2505
R21176 VSS.n4248 VSS.n2965 2.2505
R21177 VSS.n4049 VSS.n2966 2.2505
R21178 VSS.n4244 VSS.n2968 2.2505
R21179 VSS.n4243 VSS.n2969 2.2505
R21180 VSS.n4242 VSS.n2970 2.2505
R21181 VSS.n4064 VSS.n2971 2.2505
R21182 VSS.n4238 VSS.n2973 2.2505
R21183 VSS.n4237 VSS.n2974 2.2505
R21184 VSS.n4236 VSS.n2975 2.2505
R21185 VSS.n3886 VSS.n2976 2.2505
R21186 VSS.n4232 VSS.n2978 2.2505
R21187 VSS.n4231 VSS.n2979 2.2505
R21188 VSS.n4230 VSS.n2980 2.2505
R21189 VSS.n4103 VSS.n2981 2.2505
R21190 VSS.n4226 VSS.n2983 2.2505
R21191 VSS.n4225 VSS.n2984 2.2505
R21192 VSS.n4224 VSS.n2985 2.2505
R21193 VSS.n4121 VSS.n2986 2.2505
R21194 VSS.n4220 VSS.n2988 2.2505
R21195 VSS.n4219 VSS.n2989 2.2505
R21196 VSS.n4218 VSS.n2990 2.2505
R21197 VSS.n4138 VSS.n2991 2.2505
R21198 VSS.n4214 VSS.n2993 2.2505
R21199 VSS.n4213 VSS.n2994 2.2505
R21200 VSS.n4212 VSS.n2995 2.2505
R21201 VSS.n3869 VSS.n2996 2.2505
R21202 VSS.n4208 VSS.n2998 2.2505
R21203 VSS.n4207 VSS.n2999 2.2505
R21204 VSS.n4206 VSS.n3000 2.2505
R21205 VSS.n4177 VSS.n3001 2.2505
R21206 VSS.n4202 VSS.n3003 2.2505
R21207 VSS.n4201 VSS.n3004 2.2505
R21208 VSS.n4201 VSS.n3002 2.2505
R21209 VSS.n4203 VSS.n4202 2.2505
R21210 VSS.n4204 VSS.n3001 2.2505
R21211 VSS.n4206 VSS.n4205 2.2505
R21212 VSS.n4207 VSS.n2997 2.2505
R21213 VSS.n4209 VSS.n4208 2.2505
R21214 VSS.n4210 VSS.n2996 2.2505
R21215 VSS.n4212 VSS.n4211 2.2505
R21216 VSS.n4213 VSS.n2992 2.2505
R21217 VSS.n4215 VSS.n4214 2.2505
R21218 VSS.n4216 VSS.n2991 2.2505
R21219 VSS.n4218 VSS.n4217 2.2505
R21220 VSS.n4219 VSS.n2987 2.2505
R21221 VSS.n4221 VSS.n4220 2.2505
R21222 VSS.n4222 VSS.n2986 2.2505
R21223 VSS.n4224 VSS.n4223 2.2505
R21224 VSS.n4225 VSS.n2982 2.2505
R21225 VSS.n4227 VSS.n4226 2.2505
R21226 VSS.n4228 VSS.n2981 2.2505
R21227 VSS.n4230 VSS.n4229 2.2505
R21228 VSS.n4231 VSS.n2977 2.2505
R21229 VSS.n4233 VSS.n4232 2.2505
R21230 VSS.n4234 VSS.n2976 2.2505
R21231 VSS.n4236 VSS.n4235 2.2505
R21232 VSS.n4237 VSS.n2972 2.2505
R21233 VSS.n4239 VSS.n4238 2.2505
R21234 VSS.n4240 VSS.n2971 2.2505
R21235 VSS.n4242 VSS.n4241 2.2505
R21236 VSS.n4243 VSS.n2967 2.2505
R21237 VSS.n4245 VSS.n4244 2.2505
R21238 VSS.n4246 VSS.n2966 2.2505
R21239 VSS.n4248 VSS.n4247 2.2505
R21240 VSS.n4249 VSS.n2962 2.2505
R21241 VSS.n4251 VSS.n4250 2.2505
R21242 VSS.n3464 VSS.n3463 2.2505
R21243 VSS.n3461 VSS.n3460 2.2505
R21244 VSS.n3458 VSS.n3457 2.2505
R21245 VSS.n3455 VSS.n3454 2.2505
R21246 VSS.n3452 VSS.n3451 2.2505
R21247 VSS.n3449 VSS.n3448 2.2505
R21248 VSS.n3446 VSS.n2926 2.2505
R21249 VSS.n2950 VSS.n2925 2.2505
R21250 VSS.n4266 VSS.n4265 2.2505
R21251 VSS.n4263 VSS.n4262 2.2505
R21252 VSS.n4260 VSS.n4259 2.2505
R21253 VSS.n4257 VSS.n4256 2.2505
R21254 VSS.n4254 VSS.n4253 2.2505
R21255 VSS.n1796 VSS.n1523 2.2505
R21256 VSS.n2702 VSS.n1521 2.2505
R21257 VSS.n1536 VSS.n1518 2.2505
R21258 VSS.n2708 VSS.n1516 2.2505
R21259 VSS.n1540 VSS.n1513 2.2505
R21260 VSS.n2714 VSS.n1511 2.2505
R21261 VSS.n1544 VSS.n1508 2.2505
R21262 VSS.n2719 VSS.n1507 2.2505
R21263 VSS.n2721 VSS.n1505 2.2505
R21264 VSS.n2725 VSS.n1502 2.2505
R21265 VSS.n2727 VSS.n1500 2.2505
R21266 VSS.n2731 VSS.n1497 2.2505
R21267 VSS.n2733 VSS.n1495 2.2505
R21268 VSS.n2737 VSS.n1492 2.2505
R21269 VSS.n2739 VSS.n1490 2.2505
R21270 VSS.n2699 VSS.n1523 2.2505
R21271 VSS.n2702 VSS.n1519 2.2505
R21272 VSS.n2705 VSS.n1518 2.2505
R21273 VSS.n2708 VSS.n1514 2.2505
R21274 VSS.n2711 VSS.n1513 2.2505
R21275 VSS.n2714 VSS.n1509 2.2505
R21276 VSS.n2717 VSS.n1508 2.2505
R21277 VSS.n2719 VSS.n2718 2.2505
R21278 VSS.n2722 VSS.n2721 2.2505
R21279 VSS.n2725 VSS.n2724 2.2505
R21280 VSS.n2728 VSS.n2727 2.2505
R21281 VSS.n2731 VSS.n2730 2.2505
R21282 VSS.n2734 VSS.n2733 2.2505
R21283 VSS.n2737 VSS.n2736 2.2505
R21284 VSS.n2740 VSS.n2739 2.2505
R21285 VSS.n2026 VSS.n2025 2.2505
R21286 VSS.n2027 VSS.n2014 2.2505
R21287 VSS.n2181 VSS.n2006 2.2505
R21288 VSS.n2177 VSS.n1998 2.2505
R21289 VSS.n2279 VSS.n2278 2.2505
R21290 VSS.n2285 VSS.n2284 2.2505
R21291 VSS.n2307 VSS.n1959 2.2505
R21292 VSS.n1957 VSS.n1956 2.2505
R21293 VSS.n2337 VSS.n2336 2.2505
R21294 VSS.n2375 VSS.n2374 2.2505
R21295 VSS.n2385 VSS.n2384 2.2505
R21296 VSS.n2380 VSS.n1921 2.2505
R21297 VSS.n2426 VSS.n1906 2.2505
R21298 VSS.n2441 VSS.n1904 2.2505
R21299 VSS.n2473 VSS.n1892 2.2505
R21300 VSS.n2175 VSS.n2026 2.2505
R21301 VSS.n2184 VSS.n2027 2.2505
R21302 VSS.n2181 VSS.n2176 2.2505
R21303 VSS.n2178 VSS.n2177 2.2505
R21304 VSS.n2280 VSS.n2279 2.2505
R21305 VSS.n2284 VSS.n2283 2.2505
R21306 VSS.n1959 VSS.n1958 2.2505
R21307 VSS.n2334 VSS.n1957 2.2505
R21308 VSS.n2336 VSS.n2335 2.2505
R21309 VSS.n2376 VSS.n2375 2.2505
R21310 VSS.n2384 VSS.n2383 2.2505
R21311 VSS.n2381 VSS.n2380 2.2505
R21312 VSS.n1906 VSS.n1905 2.2505
R21313 VSS.n2469 VSS.n1904 2.2505
R21314 VSS.n1892 VSS.n1891 2.2505
R21315 VSS.n1525 VSS.n1524 2.2505
R21316 VSS.n2687 VSS.n2686 2.2505
R21317 VSS.n2685 VSS.n1807 2.2505
R21318 VSS.n2684 VSS.n2683 2.2505
R21319 VSS.n1809 VSS.n1808 2.2505
R21320 VSS.n2663 VSS.n2662 2.2505
R21321 VSS.n2661 VSS.n1816 2.2505
R21322 VSS.n2660 VSS.n2659 2.2505
R21323 VSS.n1818 VSS.n1817 2.2505
R21324 VSS.n2633 VSS.n2632 2.2505
R21325 VSS.n2634 VSS.n2631 2.2505
R21326 VSS.n2630 VSS.n1827 2.2505
R21327 VSS.n2629 VSS.n2628 2.2505
R21328 VSS.n1829 VSS.n1828 2.2505
R21329 VSS.n2609 VSS.n2608 2.2505
R21330 VSS.n2607 VSS.n1837 2.2505
R21331 VSS.n2606 VSS.n2605 2.2505
R21332 VSS.n1839 VSS.n1838 2.2505
R21333 VSS.n2586 VSS.n2585 2.2505
R21334 VSS.n2587 VSS.n2584 2.2505
R21335 VSS.n2583 VSS.n1854 2.2505
R21336 VSS.n2582 VSS.n2581 2.2505
R21337 VSS.n1856 VSS.n1855 2.2505
R21338 VSS.n2555 VSS.n2554 2.2505
R21339 VSS.n2556 VSS.n2553 2.2505
R21340 VSS.n2552 VSS.n1866 2.2505
R21341 VSS.n2551 VSS.n2550 2.2505
R21342 VSS.n1868 VSS.n1867 2.2505
R21343 VSS.n2531 VSS.n2530 2.2505
R21344 VSS.n2529 VSS.n1880 2.2505
R21345 VSS.n2528 VSS.n2527 2.2505
R21346 VSS.n1882 VSS.n1881 2.2505
R21347 VSS.n2509 VSS.n2508 2.2505
R21348 VSS.n2507 VSS.n1890 2.2505
R21349 VSS.n1527 VSS.n1525 2.2505
R21350 VSS.n2688 VSS.n2687 2.2505
R21351 VSS.n2675 VSS.n1807 2.2505
R21352 VSS.n2683 VSS.n2682 2.2505
R21353 VSS.n2667 VSS.n1809 2.2505
R21354 VSS.n2664 VSS.n2663 2.2505
R21355 VSS.n2652 VSS.n1816 2.2505
R21356 VSS.n2659 VSS.n2658 2.2505
R21357 VSS.n2643 VSS.n1818 2.2505
R21358 VSS.n2633 VSS.n1824 2.2505
R21359 VSS.n2635 VSS.n2634 2.2505
R21360 VSS.n2617 VSS.n1827 2.2505
R21361 VSS.n2628 VSS.n2627 2.2505
R21362 VSS.n2612 VSS.n1829 2.2505
R21363 VSS.n2610 VSS.n2609 2.2505
R21364 VSS.n1845 VSS.n1837 2.2505
R21365 VSS.n2605 VSS.n2604 2.2505
R21366 VSS.n2596 VSS.n1839 2.2505
R21367 VSS.n2586 VSS.n1851 2.2505
R21368 VSS.n2588 VSS.n2587 2.2505
R21369 VSS.n2570 VSS.n1854 2.2505
R21370 VSS.n2581 VSS.n2580 2.2505
R21371 VSS.n2565 VSS.n1856 2.2505
R21372 VSS.n2555 VSS.n1863 2.2505
R21373 VSS.n2557 VSS.n2556 2.2505
R21374 VSS.n1872 VSS.n1866 2.2505
R21375 VSS.n2550 VSS.n2549 2.2505
R21376 VSS.n2535 VSS.n1868 2.2505
R21377 VSS.n2532 VSS.n2531 2.2505
R21378 VSS.n1884 VSS.n1880 2.2505
R21379 VSS.n2527 VSS.n2526 2.2505
R21380 VSS.n2513 VSS.n1882 2.2505
R21381 VSS.n2510 VSS.n2509 2.2505
R21382 VSS.n2493 VSS.n1890 2.2505
R21383 VSS.n2074 VSS.n1441 2.2505
R21384 VSS.n2145 VSS.n2144 2.2505
R21385 VSS.n2085 VSS.n2067 2.2505
R21386 VSS.n2149 VSS.n2066 2.2505
R21387 VSS.n2150 VSS.n2065 2.2505
R21388 VSS.n2151 VSS.n2064 2.2505
R21389 VSS.n2091 VSS.n2062 2.2505
R21390 VSS.n2155 VSS.n2061 2.2505
R21391 VSS.n2156 VSS.n2060 2.2505
R21392 VSS.n2157 VSS.n2059 2.2505
R21393 VSS.n2097 VSS.n2057 2.2505
R21394 VSS.n2162 VSS.n2161 2.2505
R21395 VSS.n2054 VSS.n2029 2.2505
R21396 VSS.n2743 VSS.n1487 2.2505
R21397 VSS.n2744 VSS.n1486 2.2505
R21398 VSS.n2745 VSS.n1485 2.2505
R21399 VSS.n1627 VSS.n1483 2.2505
R21400 VSS.n2749 VSS.n1482 2.2505
R21401 VSS.n2750 VSS.n1481 2.2505
R21402 VSS.n2751 VSS.n1480 2.2505
R21403 VSS.n1606 VSS.n1478 2.2505
R21404 VSS.n2755 VSS.n1477 2.2505
R21405 VSS.n2756 VSS.n1476 2.2505
R21406 VSS.n2757 VSS.n1475 2.2505
R21407 VSS.n1585 VSS.n1471 2.2505
R21408 VSS.n2762 VSS.n2761 2.2505
R21409 VSS.n1470 VSS.n1465 2.2505
R21410 VSS.n1463 VSS.n1442 2.2505
R21411 VSS.n2743 VSS.n2742 2.2505
R21412 VSS.n2744 VSS.n1484 2.2505
R21413 VSS.n2746 VSS.n2745 2.2505
R21414 VSS.n2747 VSS.n1483 2.2505
R21415 VSS.n2749 VSS.n2748 2.2505
R21416 VSS.n2750 VSS.n1479 2.2505
R21417 VSS.n2752 VSS.n2751 2.2505
R21418 VSS.n2753 VSS.n1478 2.2505
R21419 VSS.n2755 VSS.n2754 2.2505
R21420 VSS.n2756 VSS.n1474 2.2505
R21421 VSS.n2758 VSS.n2757 2.2505
R21422 VSS.n2759 VSS.n1471 2.2505
R21423 VSS.n2761 VSS.n2760 2.2505
R21424 VSS.n1473 VSS.n1470 2.2505
R21425 VSS.n1472 VSS.n1442 2.2505
R21426 VSS.n2068 VSS.n1441 2.2505
R21427 VSS.n2146 VSS.n2145 2.2505
R21428 VSS.n2147 VSS.n2067 2.2505
R21429 VSS.n2149 VSS.n2148 2.2505
R21430 VSS.n2150 VSS.n2063 2.2505
R21431 VSS.n2152 VSS.n2151 2.2505
R21432 VSS.n2153 VSS.n2062 2.2505
R21433 VSS.n2155 VSS.n2154 2.2505
R21434 VSS.n2156 VSS.n2058 2.2505
R21435 VSS.n2158 VSS.n2157 2.2505
R21436 VSS.n2159 VSS.n2057 2.2505
R21437 VSS.n2161 VSS.n2160 2.2505
R21438 VSS.n2029 VSS.n2028 2.2505
R21439 VSS.n2802 VSS.n1445 2.2505
R21440 VSS.n2802 VSS.n1447 2.2505
R21441 VSS.n2802 VSS.n1444 2.2505
R21442 VSS.n2802 VSS.n1448 2.2505
R21443 VSS.n2802 VSS.n1443 2.2505
R21444 VSS.n2802 VSS.n2801 2.2505
R21445 VSS.n4290 VSS.n2930 2.2505
R21446 VSS.n4290 VSS.n2927 2.2505
R21447 VSS.n4028 VSS.n4027 2.2005
R21448 VSS.n4016 VSS.n4015 2.2005
R21449 VSS.n4014 VSS.n4013 2.2005
R21450 VSS.n4007 VSS.n4006 2.2005
R21451 VSS.n4005 VSS.n4004 2.2005
R21452 VSS.n3998 VSS.n3914 2.2005
R21453 VSS.n3989 VSS.n3918 2.2005
R21454 VSS.n3991 VSS.n3990 2.2005
R21455 VSS.n3987 VSS.n3986 2.2005
R21456 VSS.n3981 VSS.n3921 2.2005
R21457 VSS.n3927 VSS.n3924 2.2005
R21458 VSS.n3974 VSS.n3928 2.2005
R21459 VSS.n3969 VSS.n3968 2.2005
R21460 VSS.n3967 VSS.n3966 2.2005
R21461 VSS.n3961 VSS.n3960 2.2005
R21462 VSS.n3959 VSS.n3958 2.2005
R21463 VSS.n3953 VSS.n3952 2.2005
R21464 VSS.n3951 VSS.n3950 2.2005
R21465 VSS.n3944 VSS.n2946 2.2005
R21466 VSS.n4269 VSS.n4268 2.2005
R21467 VSS.n4271 VSS.n2944 2.2005
R21468 VSS.n4275 VSS.n2941 2.2005
R21469 VSS.n2940 VSS.n2937 2.2005
R21470 VSS.n4282 VSS.n2932 2.2005
R21471 VSS.n4288 VSS.n4287 2.2005
R21472 VSS.n3404 VSS.n2931 2.2005
R21473 VSS.n3406 VSS.n3400 2.2005
R21474 VSS.n3411 VSS.n3397 2.2005
R21475 VSS.n3396 VSS.n3394 2.2005
R21476 VSS.n3419 VSS.n3418 2.2005
R21477 VSS.n3424 VSS.n3391 2.2005
R21478 VSS.n3390 VSS.n3389 2.2005
R21479 VSS.n3431 VSS.n3386 2.2005
R21480 VSS.n3385 VSS.n3382 2.2005
R21481 VSS.n3438 VSS.n3211 2.2005
R21482 VSS.n3443 VSS.n3442 2.2005
R21483 VSS.n3377 VSS.n3210 2.2005
R21484 VSS.n3216 VSS.n3215 2.2005
R21485 VSS.n3369 VSS.n3368 2.2005
R21486 VSS.n3367 VSS.n3366 2.2005
R21487 VSS.n3360 VSS.n3359 2.2005
R21488 VSS.n3358 VSS.n3357 2.2005
R21489 VSS.n3352 VSS.n3351 2.2005
R21490 VSS.n3350 VSS.n3349 2.2005
R21491 VSS.n3343 VSS.n3226 2.2005
R21492 VSS.n3337 VSS.n3336 2.2005
R21493 VSS.n3334 VSS.n3333 2.2005
R21494 VSS.n3324 VSS.n3231 2.2005
R21495 VSS.n3326 VSS.n3325 2.2005
R21496 VSS.n3319 VSS.n3318 2.2005
R21497 VSS.n3317 VSS.n3316 2.2005
R21498 VSS.n3310 VSS.n3309 2.2005
R21499 VSS.n3308 VSS.n3307 2.2005
R21500 VSS.n3301 VSS.n3300 2.2005
R21501 VSS.n3299 VSS.n3298 2.2005
R21502 VSS.n3293 VSS.n3292 2.2005
R21503 VSS.n3291 VSS.n3290 2.2005
R21504 VSS.n3284 VSS.n3246 2.2005
R21505 VSS.n3275 VSS.n3250 2.2005
R21506 VSS.n3277 VSS.n3276 2.2005
R21507 VSS.n3270 VSS.n3269 2.2005
R21508 VSS.n3862 VSS.n3861 2.2005
R21509 VSS.n3698 VSS.n3697 2.2005
R21510 VSS.n3699 VSS.n3086 2.2005
R21511 VSS.n3702 VSS.n3701 2.2005
R21512 VSS.n3704 VSS.n3085 2.2005
R21513 VSS.n3706 VSS.n3705 2.2005
R21514 VSS.n3082 VSS.n3080 2.2005
R21515 VSS.n3718 VSS.n3717 2.2005
R21516 VSS.n3083 VSS.n3081 2.2005
R21517 VSS.n3711 VSS.n3710 2.2005
R21518 VSS.n3712 VSS.n3075 2.2005
R21519 VSS.n3727 VSS.n3074 2.2005
R21520 VSS.n3729 VSS.n3728 2.2005
R21521 VSS.n3732 VSS.n3731 2.2005
R21522 VSS.n3733 VSS.n3071 2.2005
R21523 VSS.n3736 VSS.n3735 2.2005
R21524 VSS.n3072 VSS.n3066 2.2005
R21525 VSS.n3751 VSS.n3750 2.2005
R21526 VSS.n3749 VSS.n3067 2.2005
R21527 VSS.n3748 VSS.n3747 2.2005
R21528 VSS.n3745 VSS.n3744 2.2005
R21529 VSS.n3743 VSS.n3061 2.2005
R21530 VSS.n3760 VSS.n3060 2.2005
R21531 VSS.n3762 VSS.n3761 2.2005
R21532 VSS.n3765 VSS.n3764 2.2005
R21533 VSS.n3766 VSS.n3058 2.2005
R21534 VSS.n3769 VSS.n3768 2.2005
R21535 VSS.n3049 VSS.n3047 2.2005
R21536 VSS.n3775 VSS.n3774 2.2005
R21537 VSS.n3056 VSS.n3048 2.2005
R21538 VSS.n3055 VSS.n3054 2.2005
R21539 VSS.n3052 VSS.n3051 2.2005
R21540 VSS.n3050 VSS.n3043 2.2005
R21541 VSS.n3783 VSS.n3042 2.2005
R21542 VSS.n3787 VSS.n3786 2.2005
R21543 VSS.n3784 VSS.n3040 2.2005
R21544 VSS.n3792 VSS.n3038 2.2005
R21545 VSS.n3799 VSS.n3798 2.2005
R21546 VSS.n3797 VSS.n3039 2.2005
R21547 VSS.n3795 VSS.n3794 2.2005
R21548 VSS.n3033 VSS.n3032 2.2005
R21549 VSS.n3812 VSS.n3811 2.2005
R21550 VSS.n3810 VSS.n3030 2.2005
R21551 VSS.n3818 VSS.n3817 2.2005
R21552 VSS.n3819 VSS.n3028 2.2005
R21553 VSS.n3821 VSS.n3820 2.2005
R21554 VSS.n3824 VSS.n3823 2.2005
R21555 VSS.n3825 VSS.n3026 2.2005
R21556 VSS.n3828 VSS.n3827 2.2005
R21557 VSS.n3024 VSS.n3021 2.2005
R21558 VSS.n3837 VSS.n3836 2.2005
R21559 VSS.n3835 VSS.n3023 2.2005
R21560 VSS.n3834 VSS.n3017 2.2005
R21561 VSS.n3846 VSS.n3845 2.2005
R21562 VSS.n3847 VSS.n3015 2.2005
R21563 VSS.n3850 VSS.n3849 2.2005
R21564 VSS.n3852 VSS.n3014 2.2005
R21565 VSS.n3854 VSS.n3853 2.2005
R21566 VSS.n3011 VSS.n3009 2.2005
R21567 VSS.n4194 VSS.n4193 2.2005
R21568 VSS.n3012 VSS.n3010 2.2005
R21569 VSS.n3256 VSS.n3194 2.2005
R21570 VSS.n3471 VSS.n3193 2.2005
R21571 VSS.n3473 VSS.n3472 2.2005
R21572 VSS.n3480 VSS.n3479 2.2005
R21573 VSS.n3481 VSS.n3187 2.2005
R21574 VSS.n3484 VSS.n3483 2.2005
R21575 VSS.n3486 VSS.n3185 2.2005
R21576 VSS.n3489 VSS.n3488 2.2005
R21577 VSS.n3181 VSS.n3180 2.2005
R21578 VSS.n3499 VSS.n3497 2.2005
R21579 VSS.n3176 VSS.n3175 2.2005
R21580 VSS.n3506 VSS.n3505 2.2005
R21581 VSS.n3509 VSS.n3508 2.2005
R21582 VSS.n3511 VSS.n3172 2.2005
R21583 VSS.n3514 VSS.n3513 2.2005
R21584 VSS.n3173 VSS.n3164 2.2005
R21585 VSS.n3534 VSS.n3533 2.2005
R21586 VSS.n3532 VSS.n3165 2.2005
R21587 VSS.n3168 VSS.n3167 2.2005
R21588 VSS.n3524 VSS.n3523 2.2005
R21589 VSS.n3527 VSS.n3526 2.2005
R21590 VSS.n3525 VSS.n3158 2.2005
R21591 VSS.n3542 VSS.n3541 2.2005
R21592 VSS.n3543 VSS.n3156 2.2005
R21593 VSS.n3546 VSS.n3545 2.2005
R21594 VSS.n3548 VSS.n3153 2.2005
R21595 VSS.n3560 VSS.n3559 2.2005
R21596 VSS.n3557 VSS.n3154 2.2005
R21597 VSS.n3552 VSS.n3551 2.2005
R21598 VSS.n3149 VSS.n3147 2.2005
R21599 VSS.n3572 VSS.n3571 2.2005
R21600 VSS.n3570 VSS.n3148 2.2005
R21601 VSS.n3568 VSS.n3144 2.2005
R21602 VSS.n3577 VSS.n3136 2.2005
R21603 VSS.n3580 VSS.n3579 2.2005
R21604 VSS.n3139 VSS.n3138 2.2005
R21605 VSS.n3131 VSS.n3129 2.2005
R21606 VSS.n3599 VSS.n3598 2.2005
R21607 VSS.n3132 VSS.n3130 2.2005
R21608 VSS.n3590 VSS.n3589 2.2005
R21609 VSS.n3593 VSS.n3592 2.2005
R21610 VSS.n3124 VSS.n3122 2.2005
R21611 VSS.n3607 VSS.n3606 2.2005
R21612 VSS.n3610 VSS.n3609 2.2005
R21613 VSS.n3612 VSS.n3118 2.2005
R21614 VSS.n3621 VSS.n3620 2.2005
R21615 VSS.n3618 VSS.n3119 2.2005
R21616 VSS.n3616 VSS.n3615 2.2005
R21617 VSS.n3114 VSS.n3113 2.2005
R21618 VSS.n3635 VSS.n3634 2.2005
R21619 VSS.n3633 VSS.n3111 2.2005
R21620 VSS.n3641 VSS.n3640 2.2005
R21621 VSS.n3643 VSS.n3642 2.2005
R21622 VSS.n3646 VSS.n3645 2.2005
R21623 VSS.n3647 VSS.n3106 2.2005
R21624 VSS.n3650 VSS.n3649 2.2005
R21625 VSS.n3103 VSS.n3101 2.2005
R21626 VSS.n3670 VSS.n3669 2.2005
R21627 VSS.n3653 VSS.n3102 2.2005
R21628 VSS.n3657 VSS.n3656 2.2005
R21629 VSS.n3659 VSS.n3097 2.2005
R21630 VSS.n3678 VSS.n3096 2.2005
R21631 VSS.n3681 VSS.n3680 2.2005
R21632 VSS.n3093 VSS.n3092 2.2005
R21633 VSS.n3689 VSS.n3688 2.2005
R21634 VSS.n4030 VSS.n4029 2.2005
R21635 VSS.n4039 VSS.n4038 2.2005
R21636 VSS.n4041 VSS.n4040 2.2005
R21637 VSS.n4043 VSS.n4042 2.2005
R21638 VSS.n4045 VSS.n4044 2.2005
R21639 VSS.n4046 VSS.n3895 2.2005
R21640 VSS.n4048 VSS.n4047 2.2005
R21641 VSS.n4051 VSS.n4050 2.2005
R21642 VSS.n4053 VSS.n4052 2.2005
R21643 VSS.n4055 VSS.n4054 2.2005
R21644 VSS.n4057 VSS.n4056 2.2005
R21645 VSS.n4059 VSS.n4058 2.2005
R21646 VSS.n4060 VSS.n3891 2.2005
R21647 VSS.n4063 VSS.n4062 2.2005
R21648 VSS.n4065 VSS.n3890 2.2005
R21649 VSS.n4067 VSS.n4066 2.2005
R21650 VSS.n4070 VSS.n4069 2.2005
R21651 VSS.n4068 VSS.n3888 2.2005
R21652 VSS.n4078 VSS.n4077 2.2005
R21653 VSS.n4080 VSS.n4079 2.2005
R21654 VSS.n4082 VSS.n4081 2.2005
R21655 VSS.n4084 VSS.n4083 2.2005
R21656 VSS.n4086 VSS.n4085 2.2005
R21657 VSS.n4088 VSS.n4087 2.2005
R21658 VSS.n4090 VSS.n4089 2.2005
R21659 VSS.n4092 VSS.n4091 2.2005
R21660 VSS.n4094 VSS.n4093 2.2005
R21661 VSS.n4096 VSS.n4095 2.2005
R21662 VSS.n3882 VSS.n3881 2.2005
R21663 VSS.n4102 VSS.n4101 2.2005
R21664 VSS.n4104 VSS.n3880 2.2005
R21665 VSS.n4106 VSS.n4105 2.2005
R21666 VSS.n4108 VSS.n4107 2.2005
R21667 VSS.n4110 VSS.n4109 2.2005
R21668 VSS.n4112 VSS.n4111 2.2005
R21669 VSS.n4114 VSS.n4113 2.2005
R21670 VSS.n3878 VSS.n3877 2.2005
R21671 VSS.n4120 VSS.n4119 2.2005
R21672 VSS.n4122 VSS.n3876 2.2005
R21673 VSS.n4124 VSS.n4123 2.2005
R21674 VSS.n4127 VSS.n4126 2.2005
R21675 VSS.n4129 VSS.n4128 2.2005
R21676 VSS.n4131 VSS.n4130 2.2005
R21677 VSS.n3874 VSS.n3873 2.2005
R21678 VSS.n4137 VSS.n4136 2.2005
R21679 VSS.n4139 VSS.n3872 2.2005
R21680 VSS.n4141 VSS.n4140 2.2005
R21681 VSS.n4144 VSS.n4143 2.2005
R21682 VSS.n4146 VSS.n4145 2.2005
R21683 VSS.n4149 VSS.n4148 2.2005
R21684 VSS.n4147 VSS.n3870 2.2005
R21685 VSS.n4156 VSS.n4155 2.2005
R21686 VSS.n4158 VSS.n4157 2.2005
R21687 VSS.n4160 VSS.n4159 2.2005
R21688 VSS.n4162 VSS.n4161 2.2005
R21689 VSS.n4164 VSS.n4163 2.2005
R21690 VSS.n4166 VSS.n4165 2.2005
R21691 VSS.n4168 VSS.n4167 2.2005
R21692 VSS.n4170 VSS.n4169 2.2005
R21693 VSS.n3865 VSS.n3864 2.2005
R21694 VSS.n4176 VSS.n4175 2.2005
R21695 VSS.n4178 VSS.n3863 2.2005
R21696 VSS.n4180 VSS.n4179 2.2005
R21697 VSS.n4183 VSS.n4182 2.2005
R21698 VSS.n4185 VSS.n4184 2.2005
R21699 VSS.n1528 VSS.n1526 2.2005
R21700 VSS.n1660 VSS.n1659 2.2005
R21701 VSS.n1662 VSS.n1661 2.2005
R21702 VSS.n1664 VSS.n1663 2.2005
R21703 VSS.n1665 VSS.n1560 2.2005
R21704 VSS.n1667 VSS.n1666 2.2005
R21705 VSS.n1669 VSS.n1668 2.2005
R21706 VSS.n1671 VSS.n1670 2.2005
R21707 VSS.n1673 VSS.n1672 2.2005
R21708 VSS.n1675 VSS.n1674 2.2005
R21709 VSS.n1677 VSS.n1676 2.2005
R21710 VSS.n1679 VSS.n1678 2.2005
R21711 VSS.n1681 VSS.n1680 2.2005
R21712 VSS.n1684 VSS.n1683 2.2005
R21713 VSS.n1686 VSS.n1685 2.2005
R21714 VSS.n1689 VSS.n1688 2.2005
R21715 VSS.n1687 VSS.n1554 2.2005
R21716 VSS.n1695 VSS.n1694 2.2005
R21717 VSS.n1696 VSS.n1552 2.2005
R21718 VSS.n1698 VSS.n1697 2.2005
R21719 VSS.n1701 VSS.n1700 2.2005
R21720 VSS.n1703 VSS.n1702 2.2005
R21721 VSS.n1706 VSS.n1705 2.2005
R21722 VSS.n1704 VSS.n1550 2.2005
R21723 VSS.n1712 VSS.n1711 2.2005
R21724 VSS.n1714 VSS.n1713 2.2005
R21725 VSS.n1716 VSS.n1715 2.2005
R21726 VSS.n1718 VSS.n1717 2.2005
R21727 VSS.n1720 VSS.n1719 2.2005
R21728 VSS.n1723 VSS.n1722 2.2005
R21729 VSS.n1721 VSS.n1546 2.2005
R21730 VSS.n1730 VSS.n1729 2.2005
R21731 VSS.n1732 VSS.n1731 2.2005
R21732 VSS.n1734 VSS.n1733 2.2005
R21733 VSS.n1736 VSS.n1735 2.2005
R21734 VSS.n1738 VSS.n1737 2.2005
R21735 VSS.n1740 VSS.n1739 2.2005
R21736 VSS.n1742 VSS.n1741 2.2005
R21737 VSS.n1744 VSS.n1743 2.2005
R21738 VSS.n1747 VSS.n1746 2.2005
R21739 VSS.n1749 VSS.n1748 2.2005
R21740 VSS.n1752 VSS.n1751 2.2005
R21741 VSS.n1750 VSS.n1541 2.2005
R21742 VSS.n1758 VSS.n1757 2.2005
R21743 VSS.n1759 VSS.n1539 2.2005
R21744 VSS.n1761 VSS.n1760 2.2005
R21745 VSS.n1764 VSS.n1763 2.2005
R21746 VSS.n1766 VSS.n1765 2.2005
R21747 VSS.n1769 VSS.n1768 2.2005
R21748 VSS.n1767 VSS.n1537 2.2005
R21749 VSS.n1777 VSS.n1776 2.2005
R21750 VSS.n1779 VSS.n1778 2.2005
R21751 VSS.n1781 VSS.n1780 2.2005
R21752 VSS.n1783 VSS.n1782 2.2005
R21753 VSS.n1785 VSS.n1784 2.2005
R21754 VSS.n1787 VSS.n1786 2.2005
R21755 VSS.n1790 VSS.n1789 2.2005
R21756 VSS.n1791 VSS.n1533 2.2005
R21757 VSS.n1793 VSS.n1792 2.2005
R21758 VSS.n1795 VSS.n1794 2.2005
R21759 VSS.n1798 VSS.n1797 2.2005
R21760 VSS.n2483 VSS.n1893 2.2005
R21761 VSS.n2474 VSS.n1900 2.2005
R21762 VSS.n2476 VSS.n2475 2.2005
R21763 VSS.n2448 VSS.n1903 2.2005
R21764 VSS.n2453 VSS.n2443 2.2005
R21765 VSS.n2442 VSS.n2439 2.2005
R21766 VSS.n2460 VSS.n1908 2.2005
R21767 VSS.n2465 VSS.n2464 2.2005
R21768 VSS.n2435 VSS.n1907 2.2005
R21769 VSS.n2433 VSS.n1913 2.2005
R21770 VSS.n2428 VSS.n2427 2.2005
R21771 VSS.n2425 VSS.n2424 2.2005
R21772 VSS.n2418 VSS.n2417 2.2005
R21773 VSS.n2416 VSS.n2415 2.2005
R21774 VSS.n2410 VSS.n2409 2.2005
R21775 VSS.n2408 VSS.n2407 2.2005
R21776 VSS.n2402 VSS.n2401 2.2005
R21777 VSS.n2400 VSS.n2399 2.2005
R21778 VSS.n2393 VSS.n1930 2.2005
R21779 VSS.n2387 VSS.n2386 2.2005
R21780 VSS.n1936 VSS.n1935 2.2005
R21781 VSS.n2367 VSS.n1943 2.2005
R21782 VSS.n2373 VSS.n2372 2.2005
R21783 VSS.n2361 VSS.n1941 2.2005
R21784 VSS.n2355 VSS.n2354 2.2005
R21785 VSS.n2352 VSS.n2351 2.2005
R21786 VSS.n2347 VSS.n1950 2.2005
R21787 VSS.n2338 VSS.n1953 2.2005
R21788 VSS.n2340 VSS.n2339 2.2005
R21789 VSS.n2324 VSS.n1961 2.2005
R21790 VSS.n2330 VSS.n2329 2.2005
R21791 VSS.n2317 VSS.n1960 2.2005
R21792 VSS.n2308 VSS.n1965 2.2005
R21793 VSS.n2310 VSS.n2309 2.2005
R21794 VSS.n2306 VSS.n2305 2.2005
R21795 VSS.n2299 VSS.n1968 2.2005
R21796 VSS.n1980 VSS.n1972 2.2005
R21797 VSS.n2292 VSS.n1975 2.2005
R21798 VSS.n2287 VSS.n2286 2.2005
R21799 VSS.n2270 VSS.n1978 2.2005
R21800 VSS.n1989 VSS.n1987 2.2005
R21801 VSS.n2277 VSS.n2276 2.2005
R21802 VSS.n2263 VSS.n1985 2.2005
R21803 VSS.n2257 VSS.n2256 2.2005
R21804 VSS.n2255 VSS.n2254 2.2005
R21805 VSS.n2249 VSS.n2248 2.2005
R21806 VSS.n2247 VSS.n2246 2.2005
R21807 VSS.n2242 VSS.n2241 2.2005
R21808 VSS.n2240 VSS.n2239 2.2005
R21809 VSS.n2233 VSS.n2232 2.2005
R21810 VSS.n2231 VSS.n2230 2.2005
R21811 VSS.n2223 VSS.n2222 2.2005
R21812 VSS.n2221 VSS.n2220 2.2005
R21813 VSS.n2214 VSS.n2213 2.2005
R21814 VSS.n2212 VSS.n2211 2.2005
R21815 VSS.n2206 VSS.n2205 2.2005
R21816 VSS.n2204 VSS.n2203 2.2005
R21817 VSS.n2197 VSS.n2018 2.2005
R21818 VSS.n2188 VSS.n2022 2.2005
R21819 VSS.n2190 VSS.n2189 2.2005
R21820 VSS.n2038 VSS.n2030 2.2005
R21821 VSS.n2491 VSS.n1894 2.2005
R21822 VSS.n2495 VSS.n2494 2.2005
R21823 VSS.n2496 VSS.n1889 2.2005
R21824 VSS.n2511 VSS.n1887 2.2005
R21825 VSS.n2515 VSS.n2514 2.2005
R21826 VSS.n2512 VSS.n1888 2.2005
R21827 VSS.n1885 VSS.n1883 2.2005
R21828 VSS.n2525 VSS.n2524 2.2005
R21829 VSS.n2523 VSS.n2522 2.2005
R21830 VSS.n2520 VSS.n1879 2.2005
R21831 VSS.n2533 VSS.n1876 2.2005
R21832 VSS.n2537 VSS.n2536 2.2005
R21833 VSS.n2534 VSS.n1878 2.2005
R21834 VSS.n1877 VSS.n1869 2.2005
R21835 VSS.n2548 VSS.n2547 2.2005
R21836 VSS.n2546 VSS.n1870 2.2005
R21837 VSS.n1874 VSS.n1873 2.2005
R21838 VSS.n2541 VSS.n1865 2.2005
R21839 VSS.n2558 VSS.n1864 2.2005
R21840 VSS.n2560 VSS.n2559 2.2005
R21841 VSS.n2563 VSS.n2562 2.2005
R21842 VSS.n2564 VSS.n1862 2.2005
R21843 VSS.n2567 VSS.n2566 2.2005
R21844 VSS.n1859 VSS.n1857 2.2005
R21845 VSS.n2579 VSS.n2578 2.2005
R21846 VSS.n1860 VSS.n1858 2.2005
R21847 VSS.n2572 VSS.n2571 2.2005
R21848 VSS.n2573 VSS.n1853 2.2005
R21849 VSS.n2589 VSS.n1852 2.2005
R21850 VSS.n2591 VSS.n2590 2.2005
R21851 VSS.n2594 VSS.n2593 2.2005
R21852 VSS.n2595 VSS.n1850 2.2005
R21853 VSS.n2598 VSS.n2597 2.2005
R21854 VSS.n1842 VSS.n1840 2.2005
R21855 VSS.n2603 VSS.n2602 2.2005
R21856 VSS.n1848 VSS.n1841 2.2005
R21857 VSS.n1847 VSS.n1846 2.2005
R21858 VSS.n1843 VSS.n1836 2.2005
R21859 VSS.n2611 VSS.n1835 2.2005
R21860 VSS.n2614 VSS.n2613 2.2005
R21861 VSS.n1832 VSS.n1830 2.2005
R21862 VSS.n2626 VSS.n2625 2.2005
R21863 VSS.n1833 VSS.n1831 2.2005
R21864 VSS.n2619 VSS.n2618 2.2005
R21865 VSS.n2620 VSS.n1826 2.2005
R21866 VSS.n2636 VSS.n1825 2.2005
R21867 VSS.n2638 VSS.n2637 2.2005
R21868 VSS.n2641 VSS.n2640 2.2005
R21869 VSS.n2642 VSS.n1823 2.2005
R21870 VSS.n2645 VSS.n2644 2.2005
R21871 VSS.n1821 VSS.n1819 2.2005
R21872 VSS.n2657 VSS.n2656 2.2005
R21873 VSS.n2655 VSS.n1820 2.2005
R21874 VSS.n2654 VSS.n2653 2.2005
R21875 VSS.n2650 VSS.n1815 2.2005
R21876 VSS.n2665 VSS.n1814 2.2005
R21877 VSS.n2669 VSS.n2668 2.2005
R21878 VSS.n2666 VSS.n1812 2.2005
R21879 VSS.n2674 VSS.n1810 2.2005
R21880 VSS.n2681 VSS.n2680 2.2005
R21881 VSS.n2679 VSS.n1811 2.2005
R21882 VSS.n2677 VSS.n2676 2.2005
R21883 VSS.n1806 VSS.n1805 2.2005
R21884 VSS.n2691 VSS.n2690 2.2005
R21885 VSS.n2689 VSS.n1529 2.2005
R21886 VSS.n2048 VSS.n2031 2.2005
R21887 VSS.n2055 VSS.n2052 2.2005
R21888 VSS.n2164 VSS.n2163 2.2005
R21889 VSS.n2098 VSS.n2056 2.2005
R21890 VSS.n2101 VSS.n2100 2.2005
R21891 VSS.n2103 VSS.n2102 2.2005
R21892 VSS.n2105 VSS.n2104 2.2005
R21893 VSS.n2107 VSS.n2106 2.2005
R21894 VSS.n2115 VSS.n2110 2.2005
R21895 VSS.n2117 VSS.n2116 2.2005
R21896 VSS.n2113 VSS.n2112 2.2005
R21897 VSS.n2111 VSS.n2092 2.2005
R21898 VSS.n2124 VSS.n2123 2.2005
R21899 VSS.n2126 VSS.n2125 2.2005
R21900 VSS.n2129 VSS.n2128 2.2005
R21901 VSS.n2131 VSS.n2130 2.2005
R21902 VSS.n2135 VSS.n2134 2.2005
R21903 VSS.n2133 VSS.n2132 2.2005
R21904 VSS.n2082 VSS.n2081 2.2005
R21905 VSS.n2087 VSS.n2086 2.2005
R21906 VSS.n2084 VSS.n2083 2.2005
R21907 VSS.n2071 VSS.n2069 2.2005
R21908 VSS.n2143 VSS.n2142 2.2005
R21909 VSS.n2077 VSS.n2070 2.2005
R21910 VSS.n2076 VSS.n2075 2.2005
R21911 VSS.n2072 VSS.n1449 2.2005
R21912 VSS.n2800 VSS.n2799 2.2005
R21913 VSS.n1452 VSS.n1450 2.2005
R21914 VSS.n2794 VSS.n2793 2.2005
R21915 VSS.n2792 VSS.n2791 2.2005
R21916 VSS.n2789 VSS.n2788 2.2005
R21917 VSS.n2787 VSS.n2786 2.2005
R21918 VSS.n2780 VSS.n1457 2.2005
R21919 VSS.n2782 VSS.n2781 2.2005
R21920 VSS.n2778 VSS.n2777 2.2005
R21921 VSS.n2776 VSS.n2775 2.2005
R21922 VSS.n2773 VSS.n2772 2.2005
R21923 VSS.n2771 VSS.n2770 2.2005
R21924 VSS.n2769 VSS.n2768 2.2005
R21925 VSS.n2767 VSS.n2766 2.2005
R21926 VSS.n2764 VSS.n2763 2.2005
R21927 VSS.n1580 VSS.n1469 2.2005
R21928 VSS.n1587 VSS.n1586 2.2005
R21929 VSS.n1584 VSS.n1583 2.2005
R21930 VSS.n1582 VSS.n1577 2.2005
R21931 VSS.n1594 VSS.n1593 2.2005
R21932 VSS.n1596 VSS.n1595 2.2005
R21933 VSS.n1599 VSS.n1598 2.2005
R21934 VSS.n1601 VSS.n1600 2.2005
R21935 VSS.n1609 VSS.n1608 2.2005
R21936 VSS.n1607 VSS.n1602 2.2005
R21937 VSS.n1605 VSS.n1604 2.2005
R21938 VSS.n1603 VSS.n1572 2.2005
R21939 VSS.n1617 VSS.n1616 2.2005
R21940 VSS.n1619 VSS.n1618 2.2005
R21941 VSS.n1621 VSS.n1620 2.2005
R21942 VSS.n1623 VSS.n1622 2.2005
R21943 VSS.n1630 VSS.n1629 2.2005
R21944 VSS.n1628 VSS.n1568 2.2005
R21945 VSS.n1626 VSS.n1625 2.2005
R21946 VSS.n1624 VSS.n1565 2.2005
R21947 VSS.n1641 VSS.n1640 2.2005
R21948 VSS.n1643 VSS.n1642 2.2005
R21949 VSS.n1647 VSS.n1646 2.2005
R21950 VSS.n1645 VSS.n1644 2.2005
R21951 VSS.n2907 VSS.n2906 2.15697
R21952 VSS.n736 VSS.n580 2.1255
R21953 VSS.n698 VSS.n607 2.1255
R21954 VSS.n698 VSS.n573 2.1255
R21955 VSS.n1143 VSS.n432 2.1255
R21956 VSS.n1143 VSS.n431 2.1255
R21957 VSS.n672 VSS.n671 2.11213
R21958 VSS.n1240 VSS.n365 2.0498
R21959 VSS.n1190 VSS.n419 2.04966
R21960 VSS.n736 VSS.n575 1.94252
R21961 VSS.n2909 VSS.n2908 1.9092
R21962 VSS.n1133 VSS.n1132 1.9059
R21963 VSS.n736 VSS.n735 1.86305
R21964 VSS.n831 VSS.n788 1.80449
R21965 VSS.n921 VSS.n906 1.80431
R21966 VSS.n2948 VSS.n2947 1.8005
R21967 VSS.n3935 VSS.n2949 1.8005
R21968 VSS.n4261 VSS.n2954 1.8005
R21969 VSS.n3988 VSS.n2956 1.8005
R21970 VSS.n4255 VSS.n2959 1.8005
R21971 VSS.n3462 VSS.n3198 1.8005
R21972 VSS.n3239 VSS.n3200 1.8005
R21973 VSS.n3456 VSS.n3203 1.8005
R21974 VSS.n3335 VSS.n3205 1.8005
R21975 VSS.n3450 VSS.n3208 1.8005
R21976 VSS.n3445 VSS.n3444 1.8005
R21977 VSS.n4196 VSS.n4195 1.8005
R21978 VSS.n3844 VSS.n3843 1.8005
R21979 VSS.n3839 VSS.n3838 1.8005
R21980 VSS.n3804 VSS.n3027 1.8005
R21981 VSS.n3809 VSS.n3808 1.8005
R21982 VSS.n3801 VSS.n3800 1.8005
R21983 VSS.n3053 VSS.n3044 1.8005
R21984 VSS.n3767 VSS.n3046 1.8005
R21985 VSS.n3759 VSS.n3758 1.8005
R21986 VSS.n3753 VSS.n3752 1.8005
R21987 VSS.n3077 VSS.n3073 1.8005
R21988 VSS.n3709 VSS.n3076 1.8005
R21989 VSS.n3703 VSS.n3079 1.8005
R21990 VSS.n4197 VSS.n4196 1.8005
R21991 VSS.n3843 VSS.n3842 1.8005
R21992 VSS.n3840 VSS.n3839 1.8005
R21993 VSS.n3805 VSS.n3804 1.8005
R21994 VSS.n3808 VSS.n3807 1.8005
R21995 VSS.n3802 VSS.n3801 1.8005
R21996 VSS.n3779 VSS.n3044 1.8005
R21997 VSS.n3046 VSS.n3045 1.8005
R21998 VSS.n3758 VSS.n3757 1.8005
R21999 VSS.n3754 VSS.n3753 1.8005
R22000 VSS.n3723 VSS.n3077 1.8005
R22001 VSS.n3722 VSS.n3076 1.8005
R22002 VSS.n3079 VSS.n3078 1.8005
R22003 VSS.n3693 VSS.n3089 1.8005
R22004 VSS.n3089 VSS.n3088 1.8005
R22005 VSS.n4200 VSS.n3006 1.8005
R22006 VSS.n4200 VSS.n4199 1.8005
R22007 VSS.n3462 VSS.n3196 1.8005
R22008 VSS.n3459 VSS.n3200 1.8005
R22009 VSS.n3456 VSS.n3201 1.8005
R22010 VSS.n3453 VSS.n3205 1.8005
R22011 VSS.n3450 VSS.n3206 1.8005
R22012 VSS.n3447 VSS.n3445 1.8005
R22013 VSS.n2951 VSS.n2948 1.8005
R22014 VSS.n4264 VSS.n2949 1.8005
R22015 VSS.n4261 VSS.n2952 1.8005
R22016 VSS.n4258 VSS.n2956 1.8005
R22017 VSS.n4255 VSS.n2957 1.8005
R22018 VSS.n2701 VSS.n1522 1.8005
R22019 VSS.n2703 VSS.n1520 1.8005
R22020 VSS.n2707 VSS.n1517 1.8005
R22021 VSS.n2709 VSS.n1515 1.8005
R22022 VSS.n2713 VSS.n1512 1.8005
R22023 VSS.n2715 VSS.n1510 1.8005
R22024 VSS.n2720 VSS.n1506 1.8005
R22025 VSS.n1549 VSS.n1503 1.8005
R22026 VSS.n2726 VSS.n1501 1.8005
R22027 VSS.n1553 VSS.n1498 1.8005
R22028 VSS.n2732 VSS.n1496 1.8005
R22029 VSS.n1557 VSS.n1493 1.8005
R22030 VSS.n2738 VSS.n1491 1.8005
R22031 VSS.n2701 VSS.n2700 1.8005
R22032 VSS.n2704 VSS.n2703 1.8005
R22033 VSS.n2707 VSS.n2706 1.8005
R22034 VSS.n2710 VSS.n2709 1.8005
R22035 VSS.n2713 VSS.n2712 1.8005
R22036 VSS.n2716 VSS.n2715 1.8005
R22037 VSS.n2720 VSS.n1504 1.8005
R22038 VSS.n2723 VSS.n1503 1.8005
R22039 VSS.n2726 VSS.n1499 1.8005
R22040 VSS.n2729 VSS.n1498 1.8005
R22041 VSS.n2732 VSS.n1494 1.8005
R22042 VSS.n2735 VSS.n1493 1.8005
R22043 VSS.n2738 VSS.n1489 1.8005
R22044 VSS.n2187 VSS.n2186 1.8005
R22045 VSS.n2182 VSS.n2010 1.8005
R22046 VSS.n2180 VSS.n2002 1.8005
R22047 VSS.n1994 VSS.n1984 1.8005
R22048 VSS.n1986 VSS.n1979 1.8005
R22049 VSS.n1982 VSS.n1981 1.8005
R22050 VSS.n2332 VSS.n2331 1.8005
R22051 VSS.n2353 VSS.n1940 1.8005
R22052 VSS.n1942 VSS.n1937 1.8005
R22053 VSS.n1938 VSS.n1926 1.8005
R22054 VSS.n2379 VSS.n1916 1.8005
R22055 VSS.n2467 VSS.n2466 1.8005
R22056 VSS.n2472 VSS.n2471 1.8005
R22057 VSS.n2186 VSS.n2185 1.8005
R22058 VSS.n2183 VSS.n2182 1.8005
R22059 VSS.n2180 VSS.n2179 1.8005
R22060 VSS.n1984 VSS.n1983 1.8005
R22061 VSS.n2281 VSS.n1979 1.8005
R22062 VSS.n2282 VSS.n1982 1.8005
R22063 VSS.n2333 VSS.n2332 1.8005
R22064 VSS.n1940 VSS.n1939 1.8005
R22065 VSS.n2377 VSS.n1937 1.8005
R22066 VSS.n2382 VSS.n1938 1.8005
R22067 VSS.n2379 VSS.n2378 1.8005
R22068 VSS.n2468 VSS.n2467 1.8005
R22069 VSS.n2471 VSS.n2470 1.8005
R22070 VSS.n2698 VSS.n2697 1.8005
R22071 VSS.n2697 VSS.n2696 1.8005
R22072 VSS.n1658 VSS.n1488 1.8005
R22073 VSS.n2741 VSS.n1488 1.8005
R22074 VSS.n4290 VSS.n2928 1.8005
R22075 VSS.n4290 VSS.n4289 1.8005
R22076 VSS.n95 VSS.n46 1.7762
R22077 VSS.n72 VSS.n71 1.77194
R22078 VSS.n2843 VSS.n68 1.70911
R22079 VSS.n2821 VSS.n98 1.70574
R22080 VSS.n2803 VSS.n1440 1.70453
R22081 VSS.n2901 VSS.n2900 1.704
R22082 VSS.n2903 VSS.n32 1.70222
R22083 VSS.n98 VSS.n86 1.69737
R22084 VSS.n98 VSS.n85 1.69737
R22085 VSS.n98 VSS.n97 1.6415
R22086 VSS.n735 VSS.n734 1.61453
R22087 VSS.n925 VSS.n760 1.50727
R22088 VSS.n1178 VSS.n429 1.50727
R22089 VSS.n3465 VSS.n3195 1.5005
R22090 VSS.n3268 VSS.n3195 1.5005
R22091 VSS.n4031 VSS.n2961 1.5005
R22092 VSS.n4252 VSS.n2961 1.5005
R22093 VSS.n2506 VSS.n2505 1.5005
R22094 VSS.n2505 VSS.n2504 1.5005
R22095 VSS.n2173 VSS.n2172 1.5005
R22096 VSS.n2174 VSS.n2173 1.5005
R22097 VSS.n454 VSS.n453 1.49968
R22098 VSS.n454 VSS.n452 1.49968
R22099 VSS.n1100 VSS.n446 1.49968
R22100 VSS.n1400 VSS.n1399 1.43075
R22101 VSS.n734 VSS.n575 1.4182
R22102 VSS.n1378 VSS.n155 1.41717
R22103 VSS.n747 VSS.n108 1.39698
R22104 VSS.n674 VSS.n668 1.39097
R22105 VSS.n930 VSS 1.38253
R22106 VSS.n731 VSS.n716 1.35476
R22107 VSS.n673 VSS.n669 1.3539
R22108 VSS.n2875 VSS.n2874 1.34567
R22109 VSS.n1330 VSS.n1257 1.25282
R22110 VSS VSS.n127 1.12525
R22111 VSS.n4035 VSS.n3903 1.1125
R22112 VSS.n2500 VSS.n2492 1.1125
R22113 VSS.n3663 VSS.n3658 1.10836
R22114 VSS.n1636 VSS.n1566 1.10836
R22115 VSS.n3664 VSS.n3654 1.10443
R22116 VSS.n1635 VSS.n1567 1.10443
R22117 VSS.n3687 VSS.n3686 1.10381
R22118 VSS.n1650 VSS.n1563 1.10381
R22119 VSS.n4034 VSS.n3904 1.10372
R22120 VSS.n2501 VSS.n1897 1.10372
R22121 VSS.n3668 VSS.n3667 1.10339
R22122 VSS.n1631 VSS.n1569 1.10339
R22123 VSS.n3096 VSS.n3095 1.10272
R22124 VSS.n3662 VSS.n3659 1.10272
R22125 VSS.n3665 VSS.n3653 1.10272
R22126 VSS.n1640 VSS.n1564 1.10272
R22127 VSS.n1637 VSS.n1565 1.10272
R22128 VSS.n1634 VSS.n1568 1.10272
R22129 VSS.n4038 VSS.n4037 1.10263
R22130 VSS.n4041 VSS.n3902 1.10263
R22131 VSS.n2499 VSS.n2495 1.10263
R22132 VSS.n2496 VSS.n1886 1.10263
R22133 VSS.n4192 VSS.n4191 1.1005
R22134 VSS.n3700 VSS.n3084 1.1005
R22135 VSS.n3708 VSS.n3707 1.1005
R22136 VSS.n3716 VSS.n3715 1.1005
R22137 VSS.n3714 VSS.n3713 1.1005
R22138 VSS.n3730 VSS.n3070 1.1005
R22139 VSS.n3738 VSS.n3737 1.1005
R22140 VSS.n3739 VSS.n3068 1.1005
R22141 VSS.n3740 VSS.n3069 1.1005
R22142 VSS.n3742 VSS.n3741 1.1005
R22143 VSS.n3763 VSS.n3057 1.1005
R22144 VSS.n3771 VSS.n3770 1.1005
R22145 VSS.n3773 VSS.n3772 1.1005
R22146 VSS.n3051 VSS.n3041 1.1005
R22147 VSS.n3789 VSS.n3788 1.1005
R22148 VSS.n3791 VSS.n3790 1.1005
R22149 VSS.n3796 VSS.n3031 1.1005
R22150 VSS.n3814 VSS.n3813 1.1005
R22151 VSS.n3816 VSS.n3815 1.1005
R22152 VSS.n3822 VSS.n3025 1.1005
R22153 VSS.n3830 VSS.n3829 1.1005
R22154 VSS.n3833 VSS.n3832 1.1005
R22155 VSS.n3831 VSS.n3016 1.1005
R22156 VSS.n3848 VSS.n3013 1.1005
R22157 VSS.n3856 VSS.n3855 1.1005
R22158 VSS.n3684 VSS.n3087 1.1005
R22159 VSS.n3474 VSS.n3191 1.1005
R22160 VSS.n3500 VSS.n3178 1.1005
R22161 VSS.n3555 VSS.n3554 1.1005
R22162 VSS.n3142 VSS.n3141 1.1005
R22163 VSS.n3605 VSS.n3604 1.1005
R22164 VSS.n3683 VSS.n3682 1.1005
R22165 VSS.n3661 VSS.n3660 1.1005
R22166 VSS.n3666 VSS.n3104 1.1005
R22167 VSS.n3652 VSS.n3651 1.1005
R22168 VSS.n3637 VSS.n3636 1.1005
R22169 VSS.n3603 VSS.n3123 1.1005
R22170 VSS.n3601 VSS.n3600 1.1005
R22171 VSS.n3143 VSS.n3128 1.1005
R22172 VSS.n3574 VSS.n3573 1.1005
R22173 VSS.n3556 VSS.n3146 1.1005
R22174 VSS.n3540 VSS.n3539 1.1005
R22175 VSS.n3536 VSS.n3535 1.1005
R22176 VSS.n3502 VSS.n3501 1.1005
R22177 VSS.n3478 VSS.n3477 1.1005
R22178 VSS.n3476 VSS.n3475 1.1005
R22179 VSS.n3265 VSS.n3258 1.1005
R22180 VSS.n3264 VSS.n3255 1.1005
R22181 VSS.n3257 VSS.n3192 1.1005
R22182 VSS.n3267 VSS.n3266 1.1005
R22183 VSS.n4027 VSS.n4026 1.1005
R22184 VSS.n4018 VSS.n4017 1.1005
R22185 VSS.n4016 VSS.n3909 1.1005
R22186 VSS.n4013 VSS.n4012 1.1005
R22187 VSS.n4009 VSS.n4008 1.1005
R22188 VSS.n4002 VSS.n3916 1.1005
R22189 VSS.n4004 VSS.n4003 1.1005
R22190 VSS.n4001 VSS.n3915 1.1005
R22191 VSS.n3996 VSS.n3995 1.1005
R22192 VSS.n3983 VSS.n3922 1.1005
R22193 VSS.n3982 VSS.n3981 1.1005
R22194 VSS.n3980 VSS.n3923 1.1005
R22195 VSS.n3975 VSS.n3925 1.1005
R22196 VSS.n3974 VSS.n3973 1.1005
R22197 VSS.n3972 VSS.n3926 1.1005
R22198 VSS.n3964 VSS.n3932 1.1005
R22199 VSS.n3955 VSS.n3936 1.1005
R22200 VSS.n3954 VSS.n3953 1.1005
R22201 VSS.n3938 VSS.n3937 1.1005
R22202 VSS.n3946 VSS.n3945 1.1005
R22203 VSS.n3944 VSS.n3940 1.1005
R22204 VSS.n3943 VSS.n3942 1.1005
R22205 VSS.n4270 VSS.n2943 1.1005
R22206 VSS.n4272 VSS.n4271 1.1005
R22207 VSS.n4275 VSS.n4274 1.1005
R22208 VSS.n4278 VSS.n4277 1.1005
R22209 VSS.n4281 VSS.n2936 1.1005
R22210 VSS.n4283 VSS.n4282 1.1005
R22211 VSS.n4284 VSS.n2934 1.1005
R22212 VSS.n3402 VSS.n3401 1.1005
R22213 VSS.n3410 VSS.n3409 1.1005
R22214 VSS.n3411 VSS.n3395 1.1005
R22215 VSS.n3414 VSS.n3394 1.1005
R22216 VSS.n3417 VSS.n3393 1.1005
R22217 VSS.n3422 VSS.n3392 1.1005
R22218 VSS.n3424 VSS.n3423 1.1005
R22219 VSS.n3425 VSS.n3388 1.1005
R22220 VSS.n3430 VSS.n3429 1.1005
R22221 VSS.n3437 VSS.n3381 1.1005
R22222 VSS.n3439 VSS.n3438 1.1005
R22223 VSS.n3442 VSS.n3441 1.1005
R22224 VSS.n3379 VSS.n3378 1.1005
R22225 VSS.n3375 VSS.n3374 1.1005
R22226 VSS.n3373 VSS.n3216 1.1005
R22227 VSS.n3372 VSS.n3371 1.1005
R22228 VSS.n3364 VSS.n3220 1.1005
R22229 VSS.n3354 VSS.n3223 1.1005
R22230 VSS.n3353 VSS.n3352 1.1005
R22231 VSS.n3225 VSS.n3224 1.1005
R22232 VSS.n3345 VSS.n3344 1.1005
R22233 VSS.n3343 VSS.n3228 1.1005
R22234 VSS.n3342 VSS.n3341 1.1005
R22235 VSS.n3339 VSS.n3338 1.1005
R22236 VSS.n3333 VSS.n3230 1.1005
R22237 VSS.n3330 VSS.n3231 1.1005
R22238 VSS.n3327 VSS.n3232 1.1005
R22239 VSS.n3321 VSS.n3233 1.1005
R22240 VSS.n3320 VSS.n3319 1.1005
R22241 VSS.n3235 VSS.n3234 1.1005
R22242 VSS.n3312 VSS.n3311 1.1005
R22243 VSS.n3310 VSS.n3237 1.1005
R22244 VSS.n3304 VSS.n3238 1.1005
R22245 VSS.n3303 VSS.n3240 1.1005
R22246 VSS.n3302 VSS.n3301 1.1005
R22247 VSS.n3298 VSS.n3297 1.1005
R22248 VSS.n3295 VSS.n3294 1.1005
R22249 VSS.n3288 VSS.n3248 1.1005
R22250 VSS.n3290 VSS.n3289 1.1005
R22251 VSS.n3287 VSS.n3247 1.1005
R22252 VSS.n3282 VSS.n3281 1.1005
R22253 VSS.n3272 VSS.n3252 1.1005
R22254 VSS.n3271 VSS.n3270 1.1005
R22255 VSS.n3262 VSS.n3261 1.1005
R22256 VSS.n3263 VSS.n3262 1.1005
R22257 VSS.n3260 VSS.n3255 1.1005
R22258 VSS.n3254 VSS.n3253 1.1005
R22259 VSS.n3280 VSS.n3250 1.1005
R22260 VSS.n3279 VSS.n3278 1.1005
R22261 VSS.n3277 VSS.n3251 1.1005
R22262 VSS.n3274 VSS.n3273 1.1005
R22263 VSS.n3283 VSS.n3249 1.1005
R22264 VSS.n3286 VSS.n3285 1.1005
R22265 VSS.n3245 VSS.n3244 1.1005
R22266 VSS.n3296 VSS.n3243 1.1005
R22267 VSS.n3242 VSS.n3241 1.1005
R22268 VSS.n3306 VSS.n3305 1.1005
R22269 VSS.n3313 VSS.n3236 1.1005
R22270 VSS.n3315 VSS.n3314 1.1005
R22271 VSS.n3323 VSS.n3322 1.1005
R22272 VSS.n3329 VSS.n3328 1.1005
R22273 VSS.n3332 VSS.n3331 1.1005
R22274 VSS.n3340 VSS.n3229 1.1005
R22275 VSS.n3346 VSS.n3227 1.1005
R22276 VSS.n3348 VSS.n3347 1.1005
R22277 VSS.n3356 VSS.n3355 1.1005
R22278 VSS.n3366 VSS.n3365 1.1005
R22279 VSS.n3362 VSS.n3219 1.1005
R22280 VSS.n3361 VSS.n3360 1.1005
R22281 VSS.n3222 VSS.n3221 1.1005
R22282 VSS.n3363 VSS.n3218 1.1005
R22283 VSS.n3370 VSS.n3217 1.1005
R22284 VSS.n3376 VSS.n3214 1.1005
R22285 VSS.n3380 VSS.n3212 1.1005
R22286 VSS.n3440 VSS.n3213 1.1005
R22287 VSS.n3431 VSS.n3383 1.1005
R22288 VSS.n3433 VSS.n3432 1.1005
R22289 VSS.n3434 VSS.n3382 1.1005
R22290 VSS.n3436 VSS.n3435 1.1005
R22291 VSS.n3428 VSS.n3387 1.1005
R22292 VSS.n3427 VSS.n3426 1.1005
R22293 VSS.n3421 VSS.n3420 1.1005
R22294 VSS.n3416 VSS.n3415 1.1005
R22295 VSS.n3413 VSS.n3412 1.1005
R22296 VSS.n3404 VSS.n3403 1.1005
R22297 VSS.n3405 VSS.n3399 1.1005
R22298 VSS.n3407 VSS.n3406 1.1005
R22299 VSS.n3408 VSS.n3398 1.1005
R22300 VSS.n2935 VSS.n2933 1.1005
R22301 VSS.n4286 VSS.n4285 1.1005
R22302 VSS.n4280 VSS.n4279 1.1005
R22303 VSS.n4276 VSS.n2938 1.1005
R22304 VSS.n4273 VSS.n2942 1.1005
R22305 VSS.n3941 VSS.n2945 1.1005
R22306 VSS.n3947 VSS.n3939 1.1005
R22307 VSS.n3949 VSS.n3948 1.1005
R22308 VSS.n3957 VSS.n3956 1.1005
R22309 VSS.n3966 VSS.n3965 1.1005
R22310 VSS.n3963 VSS.n3931 1.1005
R22311 VSS.n3962 VSS.n3961 1.1005
R22312 VSS.n3934 VSS.n3933 1.1005
R22313 VSS.n3930 VSS.n3929 1.1005
R22314 VSS.n3971 VSS.n3970 1.1005
R22315 VSS.n3977 VSS.n3976 1.1005
R22316 VSS.n3979 VSS.n3978 1.1005
R22317 VSS.n3986 VSS.n3985 1.1005
R22318 VSS.n3994 VSS.n3918 1.1005
R22319 VSS.n3993 VSS.n3992 1.1005
R22320 VSS.n3991 VSS.n3919 1.1005
R22321 VSS.n3984 VSS.n3920 1.1005
R22322 VSS.n3997 VSS.n3917 1.1005
R22323 VSS.n4000 VSS.n3999 1.1005
R22324 VSS.n3913 VSS.n3912 1.1005
R22325 VSS.n4010 VSS.n3911 1.1005
R22326 VSS.n4011 VSS.n3910 1.1005
R22327 VSS.n4019 VSS.n3908 1.1005
R22328 VSS.n4025 VSS.n3906 1.1005
R22329 VSS.n3907 VSS.n3905 1.1005
R22330 VSS.n4022 VSS.n4021 1.1005
R22331 VSS.n3858 VSS.n3857 1.1005
R22332 VSS.n4189 VSS.n4188 1.1005
R22333 VSS.n4190 VSS.n4189 1.1005
R22334 VSS.n4024 VSS.n3907 1.1005
R22335 VSS.n4023 VSS.n4022 1.1005
R22336 VSS.n4187 VSS.n4186 1.1005
R22337 VSS.n4181 VSS.n3859 1.1005
R22338 VSS.n4174 VSS.n4173 1.1005
R22339 VSS.n4172 VSS.n4171 1.1005
R22340 VSS.n3867 VSS.n3866 1.1005
R22341 VSS.n4152 VSS.n3868 1.1005
R22342 VSS.n4154 VSS.n4153 1.1005
R22343 VSS.n4151 VSS.n4150 1.1005
R22344 VSS.n4142 VSS.n3871 1.1005
R22345 VSS.n4135 VSS.n4134 1.1005
R22346 VSS.n4133 VSS.n4132 1.1005
R22347 VSS.n4125 VSS.n3875 1.1005
R22348 VSS.n4118 VSS.n4117 1.1005
R22349 VSS.n4116 VSS.n4115 1.1005
R22350 VSS.n4107 VSS.n3879 1.1005
R22351 VSS.n4100 VSS.n4099 1.1005
R22352 VSS.n4098 VSS.n4097 1.1005
R22353 VSS.n3884 VSS.n3883 1.1005
R22354 VSS.n4073 VSS.n3885 1.1005
R22355 VSS.n4074 VSS.n3887 1.1005
R22356 VSS.n4076 VSS.n4075 1.1005
R22357 VSS.n4072 VSS.n4071 1.1005
R22358 VSS.n4061 VSS.n3889 1.1005
R22359 VSS.n3898 VSS.n3892 1.1005
R22360 VSS.n3899 VSS.n3893 1.1005
R22361 VSS.n3900 VSS.n3894 1.1005
R22362 VSS.n3901 VSS.n3896 1.1005
R22363 VSS.n4036 VSS.n3897 1.1005
R22364 VSS.n4033 VSS.n4032 1.1005
R22365 VSS.n1800 VSS.n1799 1.1005
R22366 VSS.n1654 VSS.n1561 1.1005
R22367 VSS.n1653 VSS.n1559 1.1005
R22368 VSS.n1652 VSS.n1558 1.1005
R22369 VSS.n1651 VSS.n1556 1.1005
R22370 VSS.n1682 VSS.n1555 1.1005
R22371 VSS.n1691 VSS.n1690 1.1005
R22372 VSS.n1693 VSS.n1692 1.1005
R22373 VSS.n1699 VSS.n1551 1.1005
R22374 VSS.n1708 VSS.n1707 1.1005
R22375 VSS.n1710 VSS.n1709 1.1005
R22376 VSS.n1548 VSS.n1547 1.1005
R22377 VSS.n1725 VSS.n1724 1.1005
R22378 VSS.n1729 VSS.n1728 1.1005
R22379 VSS.n1727 VSS.n1545 1.1005
R22380 VSS.n1726 VSS.n1543 1.1005
R22381 VSS.n1745 VSS.n1542 1.1005
R22382 VSS.n1754 VSS.n1753 1.1005
R22383 VSS.n1756 VSS.n1755 1.1005
R22384 VSS.n1762 VSS.n1538 1.1005
R22385 VSS.n1771 VSS.n1770 1.1005
R22386 VSS.n1775 VSS.n1774 1.1005
R22387 VSS.n1773 VSS.n1535 1.1005
R22388 VSS.n1772 VSS.n1534 1.1005
R22389 VSS.n1788 VSS.n1532 1.1005
R22390 VSS.n1655 VSS.n1562 1.1005
R22391 VSS.n1531 VSS.n1530 1.1005
R22392 VSS.n1803 VSS.n1802 1.1005
R22393 VSS.n1802 VSS.n1801 1.1005
R22394 VSS.n2695 VSS.n2694 1.1005
R22395 VSS.n2693 VSS.n2692 1.1005
R22396 VSS.n2678 VSS.n1804 1.1005
R22397 VSS.n2673 VSS.n2672 1.1005
R22398 VSS.n2671 VSS.n2670 1.1005
R22399 VSS.n2651 VSS.n1813 1.1005
R22400 VSS.n2649 VSS.n2648 1.1005
R22401 VSS.n2647 VSS.n2646 1.1005
R22402 VSS.n2639 VSS.n1822 1.1005
R22403 VSS.n2622 VSS.n2621 1.1005
R22404 VSS.n2624 VSS.n2623 1.1005
R22405 VSS.n2616 VSS.n2615 1.1005
R22406 VSS.n1844 VSS.n1834 1.1005
R22407 VSS.n2601 VSS.n2600 1.1005
R22408 VSS.n2599 VSS.n2598 1.1005
R22409 VSS.n2592 VSS.n1849 1.1005
R22410 VSS.n2575 VSS.n2574 1.1005
R22411 VSS.n2577 VSS.n2576 1.1005
R22412 VSS.n2569 VSS.n2568 1.1005
R22413 VSS.n2561 VSS.n1861 1.1005
R22414 VSS.n2543 VSS.n2542 1.1005
R22415 VSS.n2545 VSS.n2544 1.1005
R22416 VSS.n2540 VSS.n1871 1.1005
R22417 VSS.n2539 VSS.n2538 1.1005
R22418 VSS.n2521 VSS.n1875 1.1005
R22419 VSS.n2519 VSS.n2518 1.1005
R22420 VSS.n2517 VSS.n2516 1.1005
R22421 VSS.n2498 VSS.n2497 1.1005
R22422 VSS.n2490 VSS.n1896 1.1005
R22423 VSS.n2503 VSS.n2502 1.1005
R22424 VSS.n2489 VSS.n2488 1.1005
R22425 VSS.n2486 VSS.n1896 1.1005
R22426 VSS.n2484 VSS.n2483 1.1005
R22427 VSS.n2481 VSS.n2480 1.1005
R22428 VSS.n2479 VSS.n1900 1.1005
R22429 VSS.n2476 VSS.n1901 1.1005
R22430 VSS.n2447 VSS.n2446 1.1005
R22431 VSS.n2451 VSS.n2444 1.1005
R22432 VSS.n2453 VSS.n2452 1.1005
R22433 VSS.n2454 VSS.n2440 1.1005
R22434 VSS.n2459 VSS.n2438 1.1005
R22435 VSS.n2434 VSS.n1911 1.1005
R22436 VSS.n2433 VSS.n2432 1.1005
R22437 VSS.n2431 VSS.n1912 1.1005
R22438 VSS.n2422 VSS.n1918 1.1005
R22439 VSS.n2424 VSS.n2423 1.1005
R22440 VSS.n2421 VSS.n1917 1.1005
R22441 VSS.n2413 VSS.n1923 1.1005
R22442 VSS.n2404 VSS.n1927 1.1005
R22443 VSS.n2403 VSS.n2402 1.1005
R22444 VSS.n1929 VSS.n1928 1.1005
R22445 VSS.n2395 VSS.n2394 1.1005
R22446 VSS.n2393 VSS.n1932 1.1005
R22447 VSS.n2392 VSS.n2391 1.1005
R22448 VSS.n2389 VSS.n2388 1.1005
R22449 VSS.n1935 VSS.n1934 1.1005
R22450 VSS.n2368 VSS.n2367 1.1005
R22451 VSS.n2371 VSS.n2370 1.1005
R22452 VSS.n2363 VSS.n2362 1.1005
R22453 VSS.n2361 VSS.n1946 1.1005
R22454 VSS.n2360 VSS.n2359 1.1005
R22455 VSS.n1949 VSS.n1948 1.1005
R22456 VSS.n2345 VSS.n2344 1.1005
R22457 VSS.n2343 VSS.n1953 1.1005
R22458 VSS.n2340 VSS.n1954 1.1005
R22459 VSS.n2323 VSS.n2322 1.1005
R22460 VSS.n2327 VSS.n1963 1.1005
R22461 VSS.n2329 VSS.n2328 1.1005
R22462 VSS.n2320 VSS.n1962 1.1005
R22463 VSS.n2315 VSS.n2314 1.1005
R22464 VSS.n2303 VSS.n1970 1.1005
R22465 VSS.n2305 VSS.n2304 1.1005
R22466 VSS.n2300 VSS.n2299 1.1005
R22467 VSS.n2297 VSS.n2296 1.1005
R22468 VSS.n2293 VSS.n1973 1.1005
R22469 VSS.n2292 VSS.n2291 1.1005
R22470 VSS.n2290 VSS.n1974 1.1005
R22471 VSS.n2269 VSS.n2268 1.1005
R22472 VSS.n2265 VSS.n2264 1.1005
R22473 VSS.n2263 VSS.n1990 1.1005
R22474 VSS.n2262 VSS.n2261 1.1005
R22475 VSS.n1993 VSS.n1992 1.1005
R22476 VSS.n2254 VSS.n2253 1.1005
R22477 VSS.n2252 VSS.n1995 1.1005
R22478 VSS.n1997 VSS.n1996 1.1005
R22479 VSS.n2246 VSS.n2245 1.1005
R22480 VSS.n2243 VSS.n2242 1.1005
R22481 VSS.n2238 VSS.n2237 1.1005
R22482 VSS.n2235 VSS.n2234 1.1005
R22483 VSS.n2233 VSS.n2004 1.1005
R22484 VSS.n2227 VSS.n2005 1.1005
R22485 VSS.n2225 VSS.n2224 1.1005
R22486 VSS.n2223 VSS.n2008 1.1005
R22487 VSS.n2217 VSS.n2009 1.1005
R22488 VSS.n2216 VSS.n2011 1.1005
R22489 VSS.n2215 VSS.n2214 1.1005
R22490 VSS.n2211 VSS.n2210 1.1005
R22491 VSS.n2208 VSS.n2207 1.1005
R22492 VSS.n2201 VSS.n2020 1.1005
R22493 VSS.n2203 VSS.n2202 1.1005
R22494 VSS.n2200 VSS.n2019 1.1005
R22495 VSS.n2195 VSS.n2194 1.1005
R22496 VSS.n2037 VSS.n2036 1.1005
R22497 VSS.n2039 VSS.n2038 1.1005
R22498 VSS.n2040 VSS.n2032 1.1005
R22499 VSS.n2193 VSS.n2022 1.1005
R22500 VSS.n2192 VSS.n2191 1.1005
R22501 VSS.n2190 VSS.n2023 1.1005
R22502 VSS.n2035 VSS.n2024 1.1005
R22503 VSS.n2196 VSS.n2021 1.1005
R22504 VSS.n2199 VSS.n2198 1.1005
R22505 VSS.n2017 VSS.n2016 1.1005
R22506 VSS.n2209 VSS.n2015 1.1005
R22507 VSS.n2013 VSS.n2012 1.1005
R22508 VSS.n2219 VSS.n2218 1.1005
R22509 VSS.n2226 VSS.n2007 1.1005
R22510 VSS.n2229 VSS.n2228 1.1005
R22511 VSS.n2236 VSS.n2003 1.1005
R22512 VSS.n2001 VSS.n2000 1.1005
R22513 VSS.n2244 VSS.n1999 1.1005
R22514 VSS.n2251 VSS.n2250 1.1005
R22515 VSS.n2259 VSS.n2258 1.1005
R22516 VSS.n2260 VSS.n1991 1.1005
R22517 VSS.n2266 VSS.n1988 1.1005
R22518 VSS.n2270 VSS.n2267 1.1005
R22519 VSS.n2272 VSS.n2271 1.1005
R22520 VSS.n2273 VSS.n1989 1.1005
R22521 VSS.n2275 VSS.n2274 1.1005
R22522 VSS.n1977 VSS.n1976 1.1005
R22523 VSS.n2289 VSS.n2288 1.1005
R22524 VSS.n2295 VSS.n2294 1.1005
R22525 VSS.n2298 VSS.n1971 1.1005
R22526 VSS.n2301 VSS.n1969 1.1005
R22527 VSS.n2313 VSS.n1965 1.1005
R22528 VSS.n2312 VSS.n2311 1.1005
R22529 VSS.n2310 VSS.n1966 1.1005
R22530 VSS.n2302 VSS.n1967 1.1005
R22531 VSS.n2316 VSS.n1964 1.1005
R22532 VSS.n2319 VSS.n2318 1.1005
R22533 VSS.n2326 VSS.n2325 1.1005
R22534 VSS.n2321 VSS.n1955 1.1005
R22535 VSS.n2342 VSS.n2341 1.1005
R22536 VSS.n2351 VSS.n2350 1.1005
R22537 VSS.n2349 VSS.n1951 1.1005
R22538 VSS.n2348 VSS.n2347 1.1005
R22539 VSS.n2346 VSS.n1952 1.1005
R22540 VSS.n2357 VSS.n2356 1.1005
R22541 VSS.n2358 VSS.n1947 1.1005
R22542 VSS.n2364 VSS.n1944 1.1005
R22543 VSS.n2369 VSS.n1945 1.1005
R22544 VSS.n2366 VSS.n2365 1.1005
R22545 VSS.n2390 VSS.n1933 1.1005
R22546 VSS.n2396 VSS.n1931 1.1005
R22547 VSS.n2398 VSS.n2397 1.1005
R22548 VSS.n2406 VSS.n2405 1.1005
R22549 VSS.n2415 VSS.n2414 1.1005
R22550 VSS.n2412 VSS.n1922 1.1005
R22551 VSS.n2411 VSS.n2410 1.1005
R22552 VSS.n1925 VSS.n1924 1.1005
R22553 VSS.n1920 VSS.n1919 1.1005
R22554 VSS.n2420 VSS.n2419 1.1005
R22555 VSS.n1915 VSS.n1914 1.1005
R22556 VSS.n2430 VSS.n2429 1.1005
R22557 VSS.n2436 VSS.n2435 1.1005
R22558 VSS.n2461 VSS.n2460 1.1005
R22559 VSS.n2462 VSS.n1910 1.1005
R22560 VSS.n2464 VSS.n2463 1.1005
R22561 VSS.n2437 VSS.n1909 1.1005
R22562 VSS.n2458 VSS.n2457 1.1005
R22563 VSS.n2456 VSS.n2455 1.1005
R22564 VSS.n2450 VSS.n2449 1.1005
R22565 VSS.n2445 VSS.n1902 1.1005
R22566 VSS.n2478 VSS.n2477 1.1005
R22567 VSS.n2488 VSS.n2487 1.1005
R22568 VSS.n2482 VSS.n1899 1.1005
R22569 VSS.n2485 VSS.n1895 1.1005
R22570 VSS.n2170 VSS.n2169 1.1005
R22571 VSS.n2165 VSS.n2050 1.1005
R22572 VSS.n2118 VSS.n2095 1.1005
R22573 VSS.n2795 VSS.n1453 1.1005
R22574 VSS.n1461 VSS.n1460 1.1005
R22575 VSS.n1588 VSS.n1579 1.1005
R22576 VSS.n2043 VSS.n2042 1.1005
R22577 VSS.n2045 VSS.n2033 1.1005
R22578 VSS.n2168 VSS.n2047 1.1005
R22579 VSS.n1649 VSS.n1648 1.1005
R22580 VSS.n1639 VSS.n1638 1.1005
R22581 VSS.n1633 VSS.n1632 1.1005
R22582 VSS.n1613 VSS.n1570 1.1005
R22583 VSS.n1611 VSS.n1610 1.1005
R22584 VSS.n1590 VSS.n1589 1.1005
R22585 VSS.n1466 VSS.n1462 1.1005
R22586 VSS.n1459 VSS.n1458 1.1005
R22587 VSS.n2790 VSS.n1455 1.1005
R22588 VSS.n2797 VSS.n2796 1.1005
R22589 VSS.n2141 VSS.n2140 1.1005
R22590 VSS.n2137 VSS.n2136 1.1005
R22591 VSS.n2120 VSS.n2119 1.1005
R22592 VSS.n2099 VSS.n2051 1.1005
R22593 VSS.n2167 VSS.n2166 1.1005
R22594 VSS.n2171 VSS.n2046 1.1005
R22595 VSS.n2044 VSS.n2043 1.1005
R22596 VSS.n2041 VSS.n2033 1.1005
R22597 VSS.n761 VSS.n760 1.08163
R22598 VSS.n1179 VSS.n1178 1.08163
R22599 VSS.n732 VSS.n731 1.07938
R22600 VSS.n1419 VSS.n1418 1.063
R22601 VSS.n1150 VSS 1.0355
R22602 VSS.n948 VSS.n741 0.962312
R22603 VSS.n658 VSS.n108 0.935606
R22604 VSS.n1138 VSS.n1137 0.90113
R22605 VSS VSS.n295 0.895331
R22606 VSS VSS.n164 0.895331
R22607 VSS.n1146 VSS 0.88925
R22608 VSS.n1151 VSS 0.88925
R22609 VSS.n4291 VSS.n2924 0.875
R22610 VSS.n2907 VSS 0.8695
R22611 VSS.n1100 VSS.n443 0.784892
R22612 VSS.n927 VSS.n926 0.746826
R22613 VSS.n4292 VSS.n4291 0.745657
R22614 VSS.n858 VSS.n788 0.739526
R22615 VSS.n921 VSS.n887 0.739526
R22616 VSS.n1159 VSS.n419 0.739526
R22617 VSS.n389 VSS.n365 0.739526
R22618 VSS.n3268 VSS.n3267 0.733833
R22619 VSS.n3094 VSS.n3088 0.733833
R22620 VSS.n4186 VSS.n3006 0.733833
R22621 VSS.n4032 VSS.n4031 0.733833
R22622 VSS.n2696 VSS.n2695 0.733833
R22623 VSS.n2504 VSS.n2503 0.733833
R22624 VSS.n2172 VSS.n2171 0.733833
R22625 VSS.n1658 VSS.n1657 0.733833
R22626 VSS.n846 VSS.n840 0.726116
R22627 VSS.n1252 VSS.n363 0.726116
R22628 VSS.n852 VSS.n851 0.724436
R22629 VSS.n851 VSS.n824 0.724436
R22630 VSS.n851 VSS.n821 0.724436
R22631 VSS.n787 VSS.n783 0.724436
R22632 VSS.n797 VSS.n788 0.724436
R22633 VSS.n853 VSS.n788 0.724436
R22634 VSS.n820 VSS.n788 0.724436
R22635 VSS.n823 VSS.n788 0.724436
R22636 VSS.n849 VSS.n788 0.724436
R22637 VSS.n867 VSS.n784 0.724436
R22638 VSS.n878 VSS.n780 0.724436
R22639 VSS.n921 VSS.n778 0.724436
R22640 VSS.n876 VSS.n875 0.724436
R22641 VSS.n914 VSS.n762 0.724436
R22642 VSS.n767 VSS.n762 0.724436
R22643 VSS.n765 VSS.n762 0.724436
R22644 VSS.n921 VSS.n911 0.724436
R22645 VSS.n921 VSS.n768 0.724436
R22646 VSS.n921 VSS.n766 0.724436
R22647 VSS.n921 VSS.n764 0.724436
R22648 VSS.n1174 VSS.n428 0.724436
R22649 VSS.n1170 VSS.n428 0.724436
R22650 VSS.n1168 VSS.n428 0.724436
R22651 VSS.n1173 VSS.n419 0.724436
R22652 VSS.n1169 VSS.n419 0.724436
R22653 VSS.n1167 VSS.n419 0.724436
R22654 VSS.n1220 VSS.n417 0.724436
R22655 VSS.n1222 VSS.n417 0.724436
R22656 VSS.n1223 VSS.n418 0.724436
R22657 VSS.n1219 VSS.n419 0.724436
R22658 VSS.n1233 VSS.n1232 0.724436
R22659 VSS.n1232 VSS.n411 0.724436
R22660 VSS.n378 VSS.n364 0.724436
R22661 VSS.n380 VSS.n364 0.724436
R22662 VSS.n382 VSS.n364 0.724436
R22663 VSS.n1230 VSS.n1229 0.724436
R22664 VSS.n377 VSS.n365 0.724436
R22665 VSS.n379 VSS.n365 0.724436
R22666 VSS.n381 VSS.n365 0.724436
R22667 VSS.n383 VSS.n365 0.724436
R22668 VSS.n1234 VSS.n365 0.724436
R22669 VSS.n4293 VSS.n4292 0.706573
R22670 VSS.n712 VSS.n575 0.655792
R22671 VSS.n944 VSS.n751 0.606067
R22672 VSS.n3604 VSS.n3121 0.573769
R22673 VSS.n3498 VSS.n3178 0.573769
R22674 VSS.n1581 VSS.n1579 0.573769
R22675 VSS.n2114 VSS.n2095 0.573769
R22676 VSS.n3141 VSS.n3140 0.573695
R22677 VSS.n3191 VSS.n3189 0.573695
R22678 VSS.n2774 VSS.n1461 0.573695
R22679 VSS.n2053 VSS.n2050 0.573695
R22680 VSS.n3554 VSS.n3553 0.573346
R22681 VSS.n1456 VSS.n1453 0.573346
R22682 VSS.n2784 VSS.n2783 0.573297
R22683 VSS.n3259 VSS.n3255 0.550549
R22684 VSS.n4020 VSS.n3907 0.550549
R22685 VSS.n1898 VSS.n1896 0.550549
R22686 VSS.n2034 VSS.n2033 0.550549
R22687 VSS.n2908 VSS.n2907 0.546833
R22688 VSS.n735 VSS.n584 0.53325
R22689 VSS VSS.n1144 0.517735
R22690 VSS.n1257 VSS 0.499731
R22691 VSS.n2804 VSS.n108 0.477645
R22692 VSS.n4290 VSS.n2929 0.477159
R22693 VSS.n71 VSS.n70 0.472103
R22694 VSS.n71 VSS.n69 0.472103
R22695 VSS.n71 VSS.n34 0.472103
R22696 VSS.n2901 VSS.n37 0.472103
R22697 VSS.n2901 VSS.n36 0.472103
R22698 VSS.n93 VSS.n68 0.472103
R22699 VSS.n91 VSS.n68 0.472103
R22700 VSS.n89 VSS.n68 0.472103
R22701 VSS VSS.n758 0.46028
R22702 VSS.n2901 VSS.n38 0.454928
R22703 VSS.n4291 VSS 0.398717
R22704 VSS.n987 VSS.n986 0.394692
R22705 VSS.n3603 VSS.n3125 0.39244
R22706 VSS.n3502 VSS.n3177 0.39244
R22707 VSS.n1590 VSS.n1468 0.39244
R22708 VSS.n2120 VSS.n2094 0.39244
R22709 VSS.n3578 VSS.n3128 0.389994
R22710 VSS.n3476 VSS.n3190 0.389994
R22711 VSS.n2779 VSS.n1458 0.389994
R22712 VSS.n2167 VSS.n2049 0.389994
R22713 VSS.n1149 VSS.n1148 0.389861
R22714 VSS.n1154 VSS.n1153 0.389861
R22715 VSS.n2804 VSS.n2803 0.389071
R22716 VSS.n3558 VSS.n3146 0.387191
R22717 VSS.n2798 VSS.n2797 0.387191
R22718 VSS.n1143 VSS.n433 0.385411
R22719 VSS.n3644 VSS.n3105 0.384705
R22720 VSS.n3538 VSS.n3159 0.384705
R22721 VSS.n1615 VSS.n1614 0.384705
R22722 VSS.n2139 VSS.n2078 0.384705
R22723 VSS.n3613 VSS.n3120 0.384705
R22724 VSS.n3503 VSS.n3174 0.384705
R22725 VSS.n1592 VSS.n1591 0.384705
R22726 VSS.n2122 VSS.n2121 0.384705
R22727 VSS.n3638 VSS.n3109 0.382331
R22728 VSS.n3537 VSS.n3162 0.382331
R22729 VSS.n1612 VSS.n1574 0.382331
R22730 VSS.n2138 VSS.n2088 0.382331
R22731 VSS.n3619 VSS.n3112 0.382034
R22732 VSS.n3510 VSS.n3163 0.382034
R22733 VSS.n1576 VSS.n1575 0.382034
R22734 VSS.n2090 VSS.n2089 0.382034
R22735 VSS.n3602 VSS.n3126 0.379547
R22736 VSS.n3549 VSS.n3155 0.379547
R22737 VSS.n3485 VSS.n3179 0.379547
R22738 VSS.n1467 VSS.n1464 0.379547
R22739 VSS.n1454 VSS.n1451 0.379547
R22740 VSS.n2109 VSS.n2096 0.379547
R22741 VSS.n3576 VSS.n3575 0.376968
R22742 VSS.n3575 VSS.n3145 0.376876
R22743 VSS.n3602 VSS.n3127 0.375976
R22744 VSS.n3487 VSS.n3179 0.375976
R22745 VSS.n2765 VSS.n1467 0.375976
R22746 VSS.n2109 VSS.n2108 0.375976
R22747 VSS.n3547 VSS.n3155 0.375884
R22748 VSS.n2073 VSS.n1454 0.375884
R22749 VSS.n3617 VSS.n3112 0.374982
R22750 VSS.n3512 VSS.n3163 0.374982
R22751 VSS.n1597 VSS.n1575 0.374982
R22752 VSS.n2127 VSS.n2089 0.374982
R22753 VSS.n3639 VSS.n3638 0.374889
R22754 VSS.n3537 VSS.n3161 0.374889
R22755 VSS.n1612 VSS.n1573 0.374889
R22756 VSS.n2138 VSS.n2080 0.374889
R22757 VSS.n3108 VSS.n3105 0.373984
R22758 VSS.n3538 VSS.n3160 0.373984
R22759 VSS.n1614 VSS.n1571 0.373984
R22760 VSS.n2139 VSS.n2079 0.373984
R22761 VSS.n3611 VSS.n3120 0.373891
R22762 VSS.n3504 VSS.n3503 0.373891
R22763 VSS.n1591 VSS.n1578 0.373891
R22764 VSS.n2121 VSS.n2093 0.373891
R22765 VSS.n1089 VSS.n1087 0.3701
R22766 VSS.n1075 VSS.n1074 0.3701
R22767 VSS.n1057 VSS.n1056 0.3701
R22768 VSS.n1040 VSS.n1039 0.3701
R22769 VSS.n1020 VSS.n1019 0.3701
R22770 VSS VSS.n1149 0.356592
R22771 VSS VSS.n1154 0.356592
R22772 VSS.n750 VSS.n742 0.3555
R22773 VSS.n742 VSS.n741 0.353
R22774 VSS.n1418 VSS.n155 0.344616
R22775 VSS.n2802 VSS.n1446 0.343501
R22776 VSS.n1155 VSS 0.339797
R22777 VSS.n928 VSS.n927 0.332384
R22778 VSS.n931 VSS.n930 0.332384
R22779 VSS.n950 VSS.n949 0.325527
R22780 VSS.n487 VSS.n481 0.323287
R22781 VSS.n479 VSS.n473 0.323287
R22782 VSS.n471 VSS.n465 0.323287
R22783 VSS.n1067 VSS.n1064 0.323287
R22784 VSS.n933 VSS.n759 0.300775
R22785 VSS.n1144 VSS 0.283058
R22786 VSS.n2785 VSS.n2784 0.280767
R22787 VSS.n3685 VSS.n3094 0.275034
R22788 VSS.n1657 VSS.n1656 0.275034
R22789 VSS.n1241 VSS.n1240 0.270939
R22790 VSS.n1190 VSS.n1189 0.270735
R22791 VSS VSS.n906 0.266837
R22792 VSS VSS.n831 0.266622
R22793 VSS.n951 VSS.n740 0.265372
R22794 VSS.n1096 VSS.n449 0.262114
R22795 VSS.n952 VSS.n738 0.251308
R22796 VSS.n831 VSS.n817 0.247342
R22797 VSS.n906 VSS.n905 0.247096
R22798 VSS VSS.n1190 0.245918
R22799 VSS.n1240 VSS 0.245736
R22800 VSS.n933 VSS 0.240789
R22801 VSS.n758 VSS 0.239511
R22802 VSS.n1148 VSS 0.237786
R22803 VSS.n1153 VSS 0.237786
R22804 VSS.n697 VSS.n650 0.228521
R22805 VSS.n696 VSS.n597 0.228521
R22806 VSS.n652 VSS.n649 0.228521
R22807 VSS.n661 VSS.n598 0.228521
R22808 VSS.n663 VSS.n648 0.228521
R22809 VSS.n665 VSS.n599 0.228521
R22810 VSS.n676 VSS.n600 0.228521
R22811 VSS.n678 VSS.n608 0.228521
R22812 VSS.n680 VSS.n609 0.228521
R22813 VSS.n611 VSS.n610 0.228521
R22814 VSS.n613 VSS.n586 0.228521
R22815 VSS.n612 VSS.n594 0.228521
R22816 VSS.n700 VSS.n699 0.228521
R22817 VSS.n614 VSS.n595 0.228521
R22818 VSS.n623 VSS.n615 0.228521
R22819 VSS.n646 VSS.n616 0.228521
R22820 VSS.n645 VSS.n602 0.228521
R22821 VSS.n642 VSS.n606 0.228521
R22822 VSS.n640 VSS.n603 0.228521
R22823 VSS.n638 VSS.n605 0.228521
R22824 VSS.n636 VSS.n604 0.228521
R22825 VSS.n584 VSS.n579 0.228521
R22826 VSS.n710 VSS.n578 0.228521
R22827 VSS.n711 VSS.n577 0.228521
R22828 VSS.n709 VSS.n576 0.228521
R22829 VSS.n869 VSS 0.227794
R22830 VSS.n2803 VSS 0.225507
R22831 VSS.n949 VSS.n739 0.223793
R22832 VSS.n571 VSS.n531 0.207009
R22833 VSS.n570 VSS.n524 0.207009
R22834 VSS.n567 VSS.n530 0.207009
R22835 VSS.n565 VSS.n525 0.207009
R22836 VSS.n563 VSS.n529 0.207009
R22837 VSS.n561 VSS.n527 0.207009
R22838 VSS.n559 VSS.n522 0.207009
R22839 VSS.n957 VSS.n956 0.207009
R22840 VSS.n958 VSS.n518 0.207009
R22841 VSS.n961 VSS.n960 0.207009
R22842 VSS.n517 VSS.n515 0.207009
R22843 VSS.n964 VSS.n963 0.207009
R22844 VSS.n965 VSS.n501 0.207009
R22845 VSS.n967 VSS.n502 0.207009
R22846 VSS.n969 VSS.n503 0.207009
R22847 VSS.n1000 VSS.n504 0.207009
R22848 VSS.n999 VSS.n496 0.207009
R22849 VSS.n996 VSS.n500 0.207009
R22850 VSS.n994 VSS.n497 0.207009
R22851 VSS.n992 VSS.n499 0.207009
R22852 VSS.n990 VSS.n498 0.207009
R22853 VSS.n931 VSS 0.2055
R22854 VSS.n928 VSS 0.2055
R22855 VSS.n983 VSS.n982 0.202799
R22856 VSS.n985 VSS.n984 0.202799
R22857 VSS.n984 VSS.n1 0.202799
R22858 VSS.n4294 VSS.n1 0.202799
R22859 VSS.n869 VSS 0.196087
R22860 VSS.n950 VSS.n948 0.195252
R22861 VSS.n1092 VSS.n1091 0.192746
R22862 VSS.n1102 VSS.n444 0.192746
R22863 VSS.n1070 VSS.n1068 0.192746
R22864 VSS.n1073 VSS.n1071 0.192746
R22865 VSS.n1048 VSS.n467 0.192746
R22866 VSS.n1055 VSS.n468 0.192746
R22867 VSS.n1031 VSS.n475 0.192746
R22868 VSS.n1038 VSS.n476 0.192746
R22869 VSS.n1011 VSS.n483 0.192746
R22870 VSS.n1018 VSS.n484 0.192746
R22871 VSS.n1091 VSS.n1089 0.191392
R22872 VSS.n1087 VSS.n444 0.191392
R22873 VSS.n1075 VSS.n1070 0.191392
R22874 VSS.n1074 VSS.n1073 0.191392
R22875 VSS.n1057 VSS.n467 0.191392
R22876 VSS.n1056 VSS.n1055 0.191392
R22877 VSS.n1040 VSS.n475 0.191392
R22878 VSS.n1039 VSS.n1038 0.191392
R22879 VSS.n1020 VSS.n483 0.191392
R22880 VSS.n1019 VSS.n1018 0.191392
R22881 VSS.n657 VSS.n654 0.183833
R22882 VSS.n694 VSS.n654 0.183833
R22883 VSS.n694 VSS.n655 0.183833
R22884 VSS.n690 VSS.n655 0.183833
R22885 VSS.n690 VSS.n689 0.183833
R22886 VSS.n689 VSS.n688 0.183833
R22887 VSS.n688 VSS.n667 0.183833
R22888 VSS.n683 VSS.n667 0.183833
R22889 VSS.n683 VSS.n682 0.183833
R22890 VSS.n682 VSS.n588 0.183833
R22891 VSS.n706 VSS.n588 0.183833
R22892 VSS.n706 VSS.n589 0.183833
R22893 VSS.n702 VSS.n589 0.183833
R22894 VSS.n702 VSS.n592 0.183833
R22895 VSS.n625 VSS.n592 0.183833
R22896 VSS.n626 VSS.n625 0.183833
R22897 VSS.n626 VSS.n618 0.183833
R22898 VSS.n619 VSS.n618 0.183833
R22899 VSS.n620 VSS.n619 0.183833
R22900 VSS.n621 VSS.n620 0.183833
R22901 VSS.n633 VSS.n621 0.183833
R22902 VSS.n634 VSS.n633 0.183833
R22903 VSS.n701 VSS.n593 0.183833
R22904 VSS.n624 VSS.n593 0.183833
R22905 VSS.n624 VSS.n617 0.183833
R22906 VSS.n644 VSS.n617 0.183833
R22907 VSS.n644 VSS.n643 0.183833
R22908 VSS.n643 VSS.n641 0.183833
R22909 VSS.n641 VSS.n639 0.183833
R22910 VSS.n639 VSS.n637 0.183833
R22911 VSS.n637 VSS.n635 0.183833
R22912 VSS.n656 VSS.n651 0.183833
R22913 VSS.n695 VSS.n651 0.183833
R22914 VSS.n695 VSS.n653 0.183833
R22915 VSS.n662 VSS.n653 0.183833
R22916 VSS.n664 VSS.n662 0.183833
R22917 VSS.n666 VSS.n664 0.183833
R22918 VSS.n677 VSS.n666 0.183833
R22919 VSS.n2809 VSS.n105 0.183833
R22920 VSS.n2810 VSS.n2809 0.183833
R22921 VSS.n2811 VSS.n2810 0.183833
R22922 VSS.n2811 VSS.n99 0.183833
R22923 VSS.n2819 VSS.n99 0.183833
R22924 VSS.n2820 VSS.n2819 0.183833
R22925 VSS.n2822 VSS.n78 0.183833
R22926 VSS.n2830 VSS.n78 0.183833
R22927 VSS.n2831 VSS.n2830 0.183833
R22928 VSS.n2833 VSS.n2831 0.183833
R22929 VSS.n2833 VSS.n2832 0.183833
R22930 VSS.n2842 VSS.n2841 0.183833
R22931 VSS.n2844 VSS.n62 0.183833
R22932 VSS.n2853 VSS.n62 0.183833
R22933 VSS.n2854 VSS.n2853 0.183833
R22934 VSS.n2855 VSS.n2854 0.183833
R22935 VSS.n2855 VSS.n39 0.183833
R22936 VSS.n2899 VSS.n40 0.183833
R22937 VSS.n2895 VSS.n2894 0.183833
R22938 VSS.n2894 VSS.n2893 0.183833
R22939 VSS.n2893 VSS.n47 0.183833
R22940 VSS.n2889 VSS.n47 0.183833
R22941 VSS.n2889 VSS.n2888 0.183833
R22942 VSS.n2885 VSS.n2884 0.183833
R22943 VSS.n2884 VSS.n2883 0.183833
R22944 VSS.n2883 VSS.n54 0.183833
R22945 VSS.n2879 VSS.n54 0.183833
R22946 VSS.n2879 VSS.n2878 0.183833
R22947 VSS.n2878 VSS.n14 0.183833
R22948 VSS.n759 VSS 0.180825
R22949 VSS.n1145 VSS 0.1805
R22950 VSS.n924 VSS.n761 0.174716
R22951 VSS.n1180 VSS.n1179 0.174716
R22952 VSS.n1300 VSS.n1299 0.169082
R22953 VSS.n968 VSS.n966 0.168119
R22954 VSS.n970 VSS.n968 0.168119
R22955 VSS.n970 VSS.n505 0.168119
R22956 VSS.n998 VSS.n505 0.168119
R22957 VSS.n998 VSS.n997 0.168119
R22958 VSS.n997 VSS.n995 0.168119
R22959 VSS.n995 VSS.n993 0.168119
R22960 VSS.n993 VSS.n991 0.168119
R22961 VSS.n991 VSS.n989 0.168119
R22962 VSS.n539 VSS.n532 0.168119
R22963 VSS.n569 VSS.n532 0.168119
R22964 VSS.n569 VSS.n568 0.168119
R22965 VSS.n568 VSS.n566 0.168119
R22966 VSS.n566 VSS.n564 0.168119
R22967 VSS.n564 VSS.n562 0.168119
R22968 VSS.n562 VSS.n560 0.168119
R22969 VSS VSS.n761 0.167996
R22970 VSS.n1179 VSS 0.167996
R22971 VSS.n540 VSS.n533 0.166538
R22972 VSS.n534 VSS.n533 0.166538
R22973 VSS.n535 VSS.n534 0.166538
R22974 VSS.n536 VSS.n535 0.166538
R22975 VSS.n537 VSS.n536 0.166538
R22976 VSS.n558 VSS.n537 0.166538
R22977 VSS.n558 VSS.n538 0.166538
R22978 VSS.n554 VSS.n553 0.166538
R22979 VSS.n550 VSS.n521 0.166538
R22980 VSS.n521 VSS.n514 0.166538
R22981 VSS.n514 VSS.n512 0.166538
R22982 VSS.n971 VSS.n512 0.166538
R22983 VSS.n972 VSS.n971 0.166538
R22984 VSS.n972 VSS.n506 0.166538
R22985 VSS.n507 VSS.n506 0.166538
R22986 VSS.n508 VSS.n507 0.166538
R22987 VSS.n509 VSS.n508 0.166538
R22988 VSS.n510 VSS.n509 0.166538
R22989 VSS.n988 VSS.n510 0.166538
R22990 VSS.n2821 VSS.n2820 0.1655
R22991 VSS.n1069 VSS.n1065 0.163122
R22992 VSS.n1047 VSS.n1046 0.163122
R22993 VSS.n1030 VSS.n1029 0.163122
R22994 VSS.n1010 VSS.n1009 0.163122
R22995 VSS.n1017 VSS.n1016 0.163122
R22996 VSS.n1037 VSS.n1036 0.163122
R22997 VSS.n1054 VSS.n1053 0.163122
R22998 VSS.n1072 VSS.n1061 0.163122
R22999 VSS.n1101 VSS.n445 0.163122
R23000 VSS.n949 VSS.n488 0.161915
R23001 VSS.n1060 VSS.n1059 0.158669
R23002 VSS.n1043 VSS.n1042 0.158669
R23003 VSS.n1023 VSS.n1022 0.158669
R23004 VSS.n1098 VSS.n455 0.158107
R23005 VSS.n2843 VSS.n2842 0.156333
R23006 VSS.n1072 VSS.n1062 0.154735
R23007 VSS.n1054 VSS.n469 0.154735
R23008 VSS.n1037 VSS.n477 0.154735
R23009 VSS.n1017 VSS.n485 0.154735
R23010 VSS.n2885 VSS.n32 0.1545
R23011 VSS VSS.n925 0.154142
R23012 VSS VSS.n429 0.154142
R23013 VSS.n46 VSS.n40 0.152667
R23014 VSS.n1090 VSS.n457 0.15113
R23015 VSS.n4292 VSS.n3 0.147236
R23016 VSS.n2807 VSS.n107 0.147167
R23017 VSS.n2807 VSS.n103 0.147167
R23018 VSS.n2813 VSS.n103 0.147167
R23019 VSS.n2813 VSS.n101 0.147167
R23020 VSS.n2817 VSS.n101 0.147167
R23021 VSS.n2817 VSS.n82 0.147167
R23022 VSS.n2824 VSS.n82 0.147167
R23023 VSS.n2824 VSS.n80 0.147167
R23024 VSS.n2828 VSS.n80 0.147167
R23025 VSS.n2828 VSS.n76 0.147167
R23026 VSS.n2835 VSS.n76 0.147167
R23027 VSS.n2835 VSS.n74 0.147167
R23028 VSS.n2839 VSS.n74 0.147167
R23029 VSS.n2839 VSS.n66 0.147167
R23030 VSS.n2846 VSS.n66 0.147167
R23031 VSS.n2846 VSS.n64 0.147167
R23032 VSS.n2851 VSS.n64 0.147167
R23033 VSS.n2851 VSS.n60 0.147167
R23034 VSS.n2857 VSS.n60 0.147167
R23035 VSS.n2858 VSS.n2857 0.147167
R23036 VSS.n2858 VSS.n42 0.147167
R23037 VSS.n43 VSS.n42 0.147167
R23038 VSS.n44 VSS.n43 0.147167
R23039 VSS.n2863 VSS.n44 0.147167
R23040 VSS.n2863 VSS.n48 0.147167
R23041 VSS.n49 VSS.n48 0.147167
R23042 VSS.n50 VSS.n49 0.147167
R23043 VSS.n51 VSS.n50 0.147167
R23044 VSS.n52 VSS.n51 0.147167
R23045 VSS.n2870 VSS.n52 0.147167
R23046 VSS.n2870 VSS.n55 0.147167
R23047 VSS.n56 VSS.n55 0.147167
R23048 VSS.n57 VSS.n56 0.147167
R23049 VSS.n58 VSS.n57 0.147167
R23050 VSS.n2808 VSS.n106 0.147167
R23051 VSS.n2808 VSS.n104 0.147167
R23052 VSS.n2812 VSS.n104 0.147167
R23053 VSS.n2812 VSS.n100 0.147167
R23054 VSS.n2818 VSS.n100 0.147167
R23055 VSS.n2818 VSS.n83 0.147167
R23056 VSS.n2823 VSS.n83 0.147167
R23057 VSS.n2823 VSS.n79 0.147167
R23058 VSS.n2829 VSS.n79 0.147167
R23059 VSS.n2829 VSS.n77 0.147167
R23060 VSS.n2834 VSS.n77 0.147167
R23061 VSS.n2834 VSS.n73 0.147167
R23062 VSS.n2840 VSS.n73 0.147167
R23063 VSS.n2840 VSS.n67 0.147167
R23064 VSS.n2845 VSS.n67 0.147167
R23065 VSS.n2845 VSS.n63 0.147167
R23066 VSS.n2852 VSS.n63 0.147167
R23067 VSS.n2852 VSS.n61 0.147167
R23068 VSS.n2856 VSS.n61 0.147167
R23069 VSS.n2856 VSS.n41 0.147167
R23070 VSS.n2898 VSS.n41 0.147167
R23071 VSS.n2898 VSS.n2897 0.147167
R23072 VSS.n2897 VSS.n2896 0.147167
R23073 VSS.n2896 VSS.n45 0.147167
R23074 VSS.n2892 VSS.n45 0.147167
R23075 VSS.n2892 VSS.n2891 0.147167
R23076 VSS.n2891 VSS.n2890 0.147167
R23077 VSS.n2890 VSS.n2887 0.147167
R23078 VSS.n2887 VSS.n2886 0.147167
R23079 VSS.n2886 VSS.n53 0.147167
R23080 VSS.n2882 VSS.n53 0.147167
R23081 VSS.n2882 VSS.n2881 0.147167
R23082 VSS.n2881 VSS.n2880 0.147167
R23083 VSS.n2880 VSS.n2877 0.147167
R23084 VSS.n2877 VSS.n2876 0.147167
R23085 VSS.n2900 VSS.n2899 0.145333
R23086 VSS.n2841 VSS.n72 0.141667
R23087 VSS.n1328 VSS.n1258 0.138
R23088 VSS.n1324 VSS.n1258 0.138
R23089 VSS.n1324 VSS.n1323 0.138
R23090 VSS.n1323 VSS.n1322 0.138
R23091 VSS.n1322 VSS.n1260 0.138
R23092 VSS.n1307 VSS.n1260 0.138
R23093 VSS.n1308 VSS.n1307 0.138
R23094 VSS.n1309 VSS.n1308 0.138
R23095 VSS.n1437 VSS.n112 0.138
R23096 VSS.n1433 VSS.n112 0.138
R23097 VSS.n1433 VSS.n1432 0.138
R23098 VSS.n1432 VSS.n1431 0.138
R23099 VSS.n1431 VSS.n117 0.138
R23100 VSS.n1427 VSS.n117 0.138
R23101 VSS.n1427 VSS.n1426 0.138
R23102 VSS.n1426 VSS.n1425 0.138
R23103 VSS.n1257 VSS.n1256 0.12547
R23104 VSS.n2875 VSS.n58 0.124733
R23105 VSS.n925 VSS.n924 0.12434
R23106 VSS.n1180 VSS.n429 0.12434
R23107 VSS.n447 VSS.n445 0.123672
R23108 VSS.n1069 VSS.n1066 0.123672
R23109 VSS.n1046 VSS.n464 0.123672
R23110 VSS.n1029 VSS.n472 0.123672
R23111 VSS.n1009 VSS.n480 0.123672
R23112 VSS.n1472 VSS.n1446 0.122889
R23113 VSS.n2068 VSS.n1446 0.122502
R23114 VSS.n679 VSS.n677 0.12101
R23115 VSS.n2919 VSS.n2918 0.1205
R23116 VSS.n1086 VSS.n447 0.120235
R23117 VSS.n1329 VSS.n1328 0.118364
R23118 VSS.n1425 VSS.n122 0.118364
R23119 VSS.n358 VSS 0.115394
R23120 VSS.n650 VSS.n596 0.115393
R23121 VSS.n1090 VSS.n456 0.114798
R23122 VSS.n1439 VSS.n110 0.111892
R23123 VSS.n113 VSS.n110 0.111892
R23124 VSS.n114 VSS.n113 0.111892
R23125 VSS.n115 VSS.n114 0.111892
R23126 VSS.n201 VSS.n115 0.111892
R23127 VSS.n201 VSS.n118 0.111892
R23128 VSS.n119 VSS.n118 0.111892
R23129 VSS.n120 VSS.n119 0.111892
R23130 VSS.n206 VSS.n120 0.111892
R23131 VSS.n206 VSS.n123 0.111892
R23132 VSS.n124 VSS.n123 0.111892
R23133 VSS.n125 VSS.n124 0.111892
R23134 VSS.n211 VSS.n125 0.111892
R23135 VSS.n211 VSS.n197 0.111892
R23136 VSS.n215 VSS.n197 0.111892
R23137 VSS.n215 VSS.n194 0.111892
R23138 VSS.n222 VSS.n194 0.111892
R23139 VSS.n222 VSS.n192 0.111892
R23140 VSS.n226 VSS.n192 0.111892
R23141 VSS.n226 VSS.n189 0.111892
R23142 VSS.n233 VSS.n189 0.111892
R23143 VSS.n233 VSS.n187 0.111892
R23144 VSS.n237 VSS.n187 0.111892
R23145 VSS.n237 VSS.n184 0.111892
R23146 VSS.n244 VSS.n184 0.111892
R23147 VSS.n244 VSS.n182 0.111892
R23148 VSS.n248 VSS.n182 0.111892
R23149 VSS.n248 VSS.n179 0.111892
R23150 VSS.n255 VSS.n179 0.111892
R23151 VSS.n255 VSS.n177 0.111892
R23152 VSS.n259 VSS.n177 0.111892
R23153 VSS.n259 VSS.n174 0.111892
R23154 VSS.n266 VSS.n174 0.111892
R23155 VSS.n266 VSS.n172 0.111892
R23156 VSS.n271 VSS.n172 0.111892
R23157 VSS.n271 VSS.n169 0.111892
R23158 VSS.n278 VSS.n169 0.111892
R23159 VSS.n279 VSS.n278 0.111892
R23160 VSS.n279 VSS.n160 0.111892
R23161 VSS.n161 VSS.n160 0.111892
R23162 VSS.n162 VSS.n161 0.111892
R23163 VSS.n284 VSS.n162 0.111892
R23164 VSS.n284 VSS.n165 0.111892
R23165 VSS.n1405 VSS.n165 0.111892
R23166 VSS.n1405 VSS.n1404 0.111892
R23167 VSS.n1404 VSS.n1403 0.111892
R23168 VSS.n1226 VSS 0.11175
R23169 VSS.n1088 VSS.n456 0.111609
R23170 VSS.n1398 VSS.n1397 0.1105
R23171 VSS.n1397 VSS.n291 0.1105
R23172 VSS.n293 VSS.n291 0.1105
R23173 VSS.n1266 VSS.n293 0.1105
R23174 VSS.n1266 VSS.n297 0.1105
R23175 VSS.n298 VSS.n297 0.1105
R23176 VSS.n1270 VSS.n298 0.1105
R23177 VSS.n1270 VSS.n302 0.1105
R23178 VSS.n303 VSS.n302 0.1105
R23179 VSS.n304 VSS.n303 0.1105
R23180 VSS.n1275 VSS.n304 0.1105
R23181 VSS.n1275 VSS.n332 0.1105
R23182 VSS.n333 VSS.n332 0.1105
R23183 VSS.n334 VSS.n333 0.1105
R23184 VSS.n335 VSS.n334 0.1105
R23185 VSS.n336 VSS.n335 0.1105
R23186 VSS.n337 VSS.n336 0.1105
R23187 VSS.n338 VSS.n337 0.1105
R23188 VSS.n339 VSS.n338 0.1105
R23189 VSS.n340 VSS.n339 0.1105
R23190 VSS.n341 VSS.n340 0.1105
R23191 VSS.n342 VSS.n341 0.1105
R23192 VSS.n343 VSS.n342 0.1105
R23193 VSS.n344 VSS.n343 0.1105
R23194 VSS.n345 VSS.n344 0.1105
R23195 VSS.n346 VSS.n345 0.1105
R23196 VSS.n347 VSS.n346 0.1105
R23197 VSS.n348 VSS.n347 0.1105
R23198 VSS.n349 VSS.n348 0.1105
R23199 VSS.n350 VSS.n349 0.1105
R23200 VSS.n351 VSS.n350 0.1105
R23201 VSS.n352 VSS.n351 0.1105
R23202 VSS.n353 VSS.n352 0.1105
R23203 VSS.n354 VSS.n353 0.1105
R23204 VSS.n1396 VSS.n1395 0.1105
R23205 VSS.n1395 VSS.n1394 0.1105
R23206 VSS.n1394 VSS.n294 0.1105
R23207 VSS.n1390 VSS.n294 0.1105
R23208 VSS.n1390 VSS.n1389 0.1105
R23209 VSS.n1389 VSS.n299 0.1105
R23210 VSS.n1383 VSS.n299 0.1105
R23211 VSS.n1383 VSS.n1382 0.1105
R23212 VSS.n1382 VSS.n1381 0.1105
R23213 VSS.n1381 VSS.n305 0.1105
R23214 VSS.n1375 VSS.n305 0.1105
R23215 VSS.n1375 VSS.n1374 0.1105
R23216 VSS.n1374 VSS.n1372 0.1105
R23217 VSS.n1372 VSS.n1370 0.1105
R23218 VSS.n1370 VSS.n1368 0.1105
R23219 VSS.n1368 VSS.n1366 0.1105
R23220 VSS.n1366 VSS.n1364 0.1105
R23221 VSS.n1364 VSS.n1362 0.1105
R23222 VSS.n1362 VSS.n1360 0.1105
R23223 VSS.n1360 VSS.n1358 0.1105
R23224 VSS.n1358 VSS.n1356 0.1105
R23225 VSS.n1356 VSS.n1354 0.1105
R23226 VSS.n1354 VSS.n1352 0.1105
R23227 VSS.n1352 VSS.n1350 0.1105
R23228 VSS.n1350 VSS.n1348 0.1105
R23229 VSS.n1348 VSS.n1346 0.1105
R23230 VSS.n1346 VSS.n1344 0.1105
R23231 VSS.n1344 VSS.n1342 0.1105
R23232 VSS.n1342 VSS.n1340 0.1105
R23233 VSS.n1340 VSS.n1338 0.1105
R23234 VSS.n1338 VSS.n1336 0.1105
R23235 VSS.n1336 VSS.n1334 0.1105
R23236 VSS.n1334 VSS.n1332 0.1105
R23237 VSS.n1332 VSS.n355 0.1105
R23238 VSS.n1327 VSS.n355 0.1105
R23239 VSS.n1327 VSS.n1326 0.1105
R23240 VSS.n1326 VSS.n1325 0.1105
R23241 VSS.n1325 VSS.n1259 0.1105
R23242 VSS.n1321 VSS.n1259 0.1105
R23243 VSS.n1321 VSS.n1261 0.1105
R23244 VSS.n1302 VSS.n1261 0.1105
R23245 VSS.n1303 VSS.n1302 0.1105
R23246 VSS.n1304 VSS.n1303 0.1105
R23247 VSS.n1306 VSS.n1304 0.1105
R23248 VSS.n1320 VSS.n1262 0.1105
R23249 VSS.n1320 VSS.n1263 0.1105
R23250 VSS.n1316 VSS.n1263 0.1105
R23251 VSS.n1316 VSS.n1315 0.1105
R23252 VSS.n1315 VSS.n1314 0.1105
R23253 VSS.n1314 VSS.n1305 0.1105
R23254 VSS.n1436 VSS.n111 0.1105
R23255 VSS.n1436 VSS.n1435 0.1105
R23256 VSS.n1435 VSS.n1434 0.1105
R23257 VSS.n1434 VSS.n116 0.1105
R23258 VSS.n1430 VSS.n116 0.1105
R23259 VSS.n1430 VSS.n1429 0.1105
R23260 VSS.n1429 VSS.n1428 0.1105
R23261 VSS.n1428 VSS.n121 0.1105
R23262 VSS.n1424 VSS.n121 0.1105
R23263 VSS.n1424 VSS.n1423 0.1105
R23264 VSS.n1423 VSS.n1422 0.1105
R23265 VSS.n1422 VSS.n126 0.1105
R23266 VSS.n196 VSS.n126 0.1105
R23267 VSS.n217 VSS.n196 0.1105
R23268 VSS.n219 VSS.n217 0.1105
R23269 VSS.n221 VSS.n219 0.1105
R23270 VSS.n221 VSS.n191 0.1105
R23271 VSS.n228 VSS.n191 0.1105
R23272 VSS.n230 VSS.n228 0.1105
R23273 VSS.n232 VSS.n230 0.1105
R23274 VSS.n232 VSS.n186 0.1105
R23275 VSS.n239 VSS.n186 0.1105
R23276 VSS.n241 VSS.n239 0.1105
R23277 VSS.n243 VSS.n241 0.1105
R23278 VSS.n243 VSS.n181 0.1105
R23279 VSS.n250 VSS.n181 0.1105
R23280 VSS.n252 VSS.n250 0.1105
R23281 VSS.n254 VSS.n252 0.1105
R23282 VSS.n254 VSS.n176 0.1105
R23283 VSS.n261 VSS.n176 0.1105
R23284 VSS.n263 VSS.n261 0.1105
R23285 VSS.n265 VSS.n263 0.1105
R23286 VSS.n265 VSS.n171 0.1105
R23287 VSS.n273 VSS.n171 0.1105
R23288 VSS.n275 VSS.n273 0.1105
R23289 VSS.n277 VSS.n275 0.1105
R23290 VSS.n277 VSS.n159 0.1105
R23291 VSS.n1414 VSS.n159 0.1105
R23292 VSS.n1414 VSS.n1413 0.1105
R23293 VSS.n1413 VSS.n1411 0.1105
R23294 VSS.n1411 VSS.n163 0.1105
R23295 VSS.n1407 VSS.n163 0.1105
R23296 VSS.n1407 VSS.n1406 0.1105
R23297 VSS.n1406 VSS.n167 0.1105
R23298 VSS.n2908 VSS.n14 0.108667
R23299 VSS VSS.n844 0.104833
R23300 VSS.n531 VSS.n523 0.104666
R23301 VSS.n4295 VSS.n0 0.102427
R23302 VSS.n982 VSS.n0 0.0996547
R23303 VSS.n983 VSS.n981 0.0996547
R23304 VSS.n3446 VSS.n2929 0.0982363
R23305 VSS.n2950 VSS.n2929 0.0974074
R23306 VSS.n2923 VSS.n5 0.0965
R23307 VSS.n2917 VSS.n6 0.0965
R23308 VSS.n2922 VSS.n6 0.0965
R23309 VSS VSS.n674 0.0949503
R23310 VSS.n1066 VSS.n455 0.0927349
R23311 VSS.n1059 VSS.n464 0.0927349
R23312 VSS.n1042 VSS.n472 0.0927349
R23313 VSS.n1022 VSS.n480 0.0927349
R23314 VSS.n722 VSS.n720 0.0842132
R23315 VSS.n727 VSS.n715 0.0842132
R23316 VSS.n723 VSS.n719 0.0834044
R23317 VSS.n538 VSS.n519 0.0832601
R23318 VSS.n553 VSS.n520 0.0832601
R23319 VSS.n550 VSS.n520 0.0832601
R23320 VSS.n554 VSS.n519 0.0832601
R23321 VSS.n541 VSS.n540 0.0830423
R23322 VSS.n1132 VSS.n105 0.083
R23323 VSS.n728 VSS.n726 0.0805735
R23324 VSS.n357 VSS 0.0805495
R23325 VSS.n844 VSS 0.0802977
R23326 VSS.n560 VSS.n513 0.0784429
R23327 VSS.n1311 VSS 0.0775
R23328 VSS.n1402 VSS 0.0775
R23329 VSS.n865 VSS 0.0684471
R23330 VSS.n779 VSS 0.0684471
R23331 VSS.n843 VSS.n835 0.068
R23332 VSS.n924 VSS.n923 0.068
R23333 VSS.n701 VSS.n587 0.0674674
R23334 VSS VSS.n1211 0.0649962
R23335 VSS VSS.n412 0.0649962
R23336 VSS.n1067 VSS.n1062 0.06234
R23337 VSS.n469 VSS.n465 0.06234
R23338 VSS.n477 VSS.n473 0.06234
R23339 VSS.n485 VSS.n481 0.06234
R23340 VSS.n2806 VSS.n2805 0.0616111
R23341 VSS.n2806 VSS.n102 0.0616111
R23342 VSS.n2814 VSS.n102 0.0616111
R23343 VSS.n2815 VSS.n2814 0.0616111
R23344 VSS.n2816 VSS.n2815 0.0616111
R23345 VSS.n2816 VSS.n81 0.0616111
R23346 VSS.n2825 VSS.n81 0.0616111
R23347 VSS.n2826 VSS.n2825 0.0616111
R23348 VSS.n2827 VSS.n2826 0.0616111
R23349 VSS.n2827 VSS.n75 0.0616111
R23350 VSS.n2836 VSS.n75 0.0616111
R23351 VSS.n2837 VSS.n2836 0.0616111
R23352 VSS.n2838 VSS.n2837 0.0616111
R23353 VSS.n2838 VSS.n65 0.0616111
R23354 VSS.n2847 VSS.n65 0.0616111
R23355 VSS.n2848 VSS.n2847 0.0616111
R23356 VSS.n2850 VSS.n2848 0.0616111
R23357 VSS.n2850 VSS.n2849 0.0616111
R23358 VSS.n2849 VSS.n59 0.0616111
R23359 VSS.n2859 VSS.n59 0.0616111
R23360 VSS.n2860 VSS.n2859 0.0616111
R23361 VSS.n2861 VSS.n2860 0.0616111
R23362 VSS.n2862 VSS.n2861 0.0616111
R23363 VSS.n2864 VSS.n2862 0.0616111
R23364 VSS.n2865 VSS.n2864 0.0616111
R23365 VSS.n2866 VSS.n2865 0.0616111
R23366 VSS.n2867 VSS.n2866 0.0616111
R23367 VSS.n2868 VSS.n2867 0.0616111
R23368 VSS.n2869 VSS.n2868 0.0616111
R23369 VSS.n2871 VSS.n2869 0.0616111
R23370 VSS.n2872 VSS.n2871 0.0616111
R23371 VSS.n2873 VSS.n2872 0.0616111
R23372 VSS.n2874 VSS.n2873 0.0616111
R23373 VSS.n834 VSS.n822 0.0613943
R23374 VSS.n826 VSS.n825 0.0613943
R23375 VSS.n830 VSS.n829 0.0613943
R23376 VSS.n866 VSS.n786 0.0613943
R23377 VSS.n832 VSS.n830 0.0613943
R23378 VSS.n829 VSS.n826 0.0613943
R23379 VSS.n825 VSS.n822 0.0613943
R23380 VSS.n866 VSS.n865 0.0613943
R23381 VSS.n922 VSS.n763 0.0613943
R23382 VSS.n920 VSS.n919 0.0613943
R23383 VSS.n918 VSS.n917 0.0613943
R23384 VSS.n874 VSS.n781 0.0613943
R23385 VSS.n874 VSS.n779 0.0613943
R23386 VSS.n917 VSS.n913 0.0613943
R23387 VSS.n919 VSS.n918 0.0613943
R23388 VSS.n920 VSS.n763 0.0613943
R23389 VSS.n1188 VSS.n1187 0.0613943
R23390 VSS.n1186 VSS.n1185 0.0613943
R23391 VSS.n1184 VSS.n1183 0.0613943
R23392 VSS.n1183 VSS.n1182 0.0613943
R23393 VSS.n1185 VSS.n1184 0.0613943
R23394 VSS.n1187 VSS.n1186 0.0613943
R23395 VSS.n1243 VSS.n1242 0.0613943
R23396 VSS.n1245 VSS.n1244 0.0613943
R23397 VSS.n1247 VSS.n1246 0.0613943
R23398 VSS.n1248 VSS.n1247 0.0613943
R23399 VSS.n1246 VSS.n1245 0.0613943
R23400 VSS.n1244 VSS.n1243 0.0613943
R23401 VSS.n1212 VSS 0.0609472
R23402 VSS.n415 VSS 0.0609472
R23403 VSS.n2920 VSS.n2919 0.060789
R23404 VSS.n2921 VSS.n2920 0.060789
R23405 VSS VSS.n932 0.0605
R23406 VSS VSS.n929 0.0605
R23407 VSS.n2921 VSS 0.0605
R23408 VSS.n749 VSS.n743 0.0597227
R23409 VSS.n744 VSS.n743 0.0593057
R23410 VSS VSS.n2802 0.057347
R23411 VSS.n295 VSS.n292 0.0565855
R23412 VSS.n166 VSS.n164 0.0561031
R23413 VSS.n1311 VSS.n1310 0.0560829
R23414 VSS.n1402 VSS.n1401 0.0560829
R23415 VSS.n1312 VSS.n1305 0.0555643
R23416 VSS.n1310 VSS.n1306 0.055254
R23417 VSS.n1396 VSS.n290 0.055254
R23418 VSS.n1401 VSS.n167 0.055254
R23419 VSS.n1438 VSS.n111 0.055254
R23420 VSS.n1226 VSS 0.054882
R23421 VSS.n863 VSS 0.0534472
R23422 VSS VSS.n880 0.0534472
R23423 VSS VSS.n4290 0.0533417
R23424 VSS.n817 VSS.n816 0.053
R23425 VSS.n810 VSS.n791 0.053
R23426 VSS.n812 VSS.n811 0.053
R23427 VSS.n804 VSS.n793 0.053
R23428 VSS.n806 VSS.n805 0.053
R23429 VSS.n799 VSS.n795 0.053
R23430 VSS.n800 VSS.n789 0.053
R23431 VSS.n905 VSS.n771 0.053
R23432 VSS.n890 VSS.n885 0.053
R23433 VSS.n901 VSS.n773 0.053
R23434 VSS.n892 VSS.n883 0.053
R23435 VSS.n899 VSS.n775 0.053
R23436 VSS.n894 VSS.n881 0.053
R23437 VSS.n897 VSS.n777 0.053
R23438 VSS.n1216 VSS.n1214 0.053
R23439 VSS.n1215 VSS.n422 0.053
R23440 VSS.n1207 VSS.n1205 0.053
R23441 VSS.n1206 VSS.n424 0.053
R23442 VSS.n1201 VSS.n1199 0.053
R23443 VSS.n1200 VSS.n426 0.053
R23444 VSS.n1195 VSS.n1193 0.053
R23445 VSS.n1194 VSS.n1192 0.053
R23446 VSS.n413 VSS.n409 0.053
R23447 VSS.n408 VSS.n368 0.053
R23448 VSS.n404 VSS.n402 0.053
R23449 VSS.n403 VSS.n370 0.053
R23450 VSS.n398 VSS.n396 0.053
R23451 VSS.n397 VSS.n372 0.053
R23452 VSS.n392 VSS.n391 0.053
R23453 VSS.n1238 VSS.n366 0.053
R23454 VSS.n1257 VSS 0.0520042
R23455 VSS.n1409 VSS.n1408 0.0487456
R23456 VSS.n1393 VSS.n1392 0.0487456
R23457 VSS.n1392 VSS.n1391 0.0487456
R23458 VSS.n1384 VSS.n301 0.0487456
R23459 VSS.n5 VSS.n4 0.0487454
R23460 VSS.n543 VSS.n542 0.0487192
R23461 VSS.n544 VSS.n543 0.0487192
R23462 VSS.n545 VSS.n544 0.0487192
R23463 VSS.n546 VSS.n545 0.0487192
R23464 VSS.n557 VSS.n546 0.0487192
R23465 VSS.n557 VSS.n556 0.0487192
R23466 VSS.n556 VSS.n555 0.0487192
R23467 VSS.n555 VSS.n552 0.0487192
R23468 VSS.n552 VSS.n551 0.0487192
R23469 VSS.n551 VSS.n549 0.0487192
R23470 VSS.n549 VSS.n548 0.0487192
R23471 VSS.n548 VSS.n547 0.0487192
R23472 VSS.n547 VSS.n511 0.0487192
R23473 VSS.n973 VSS.n511 0.0487192
R23474 VSS.n974 VSS.n973 0.0487192
R23475 VSS.n975 VSS.n974 0.0487192
R23476 VSS.n976 VSS.n975 0.0487192
R23477 VSS.n977 VSS.n976 0.0487192
R23478 VSS.n978 VSS.n977 0.0487192
R23479 VSS.n987 VSS.n978 0.0487192
R23480 VSS.n986 VSS.n979 0.0487192
R23481 VSS.n979 VSS.n2 0.0487192
R23482 VSS.n4293 VSS.n2 0.0487192
R23483 VSS.n842 VSS 0.048535
R23484 VSS VSS.n362 0.048535
R23485 VSS.n1097 VSS.n1096 0.0477982
R23486 VSS.n966 VSS.n513 0.0474333
R23487 VSS.n926 VSS 0.0462933
R23488 VSS.n1155 VSS 0.0462933
R23489 VSS.n251 VSS.n131 0.0458509
R23490 VSS.n253 VSS.n139 0.0458509
R23491 VSS.n1365 VSS.n310 0.0458509
R23492 VSS.n1363 VSS.n328 0.0458509
R23493 VSS VSS.n359 0.0457384
R23494 VSS.n931 VSS 0.0457336
R23495 VSS.n928 VSS 0.0457336
R23496 VSS.n249 VSS.n141 0.0439211
R23497 VSS.n175 VSS.n132 0.0439211
R23498 VSS VSS.n1409 0.0439211
R23499 VSS.n1367 VSS.n330 0.0439211
R23500 VSS.n1361 VSS.n311 0.0439211
R23501 VSS.n2832 VSS.n72 0.0426667
R23502 VSS.n180 VSS.n130 0.0419912
R23503 VSS.n1359 VSS.n325 0.0419912
R23504 VSS.n260 VSS.n138 0.0419912
R23505 VSS VSS.n158 0.0419912
R23506 VSS.n1369 VSS.n309 0.0419912
R23507 VSS.n1086 VSS.n449 0.04175
R23508 VSS.n681 VSS.n679 0.041053
R23509 VSS.n681 VSS.n585 0.041053
R23510 VSS.n707 VSS.n587 0.041053
R23511 VSS.n2948 VSS.n2925 0.0405
R23512 VSS.n4266 VSS.n2948 0.0405
R23513 VSS.n4266 VSS.n2949 0.0405
R23514 VSS.n4262 VSS.n2949 0.0405
R23515 VSS.n4262 VSS.n4261 0.0405
R23516 VSS.n4261 VSS.n4260 0.0405
R23517 VSS.n4260 VSS.n2956 0.0405
R23518 VSS.n4256 VSS.n2956 0.0405
R23519 VSS.n4256 VSS.n4255 0.0405
R23520 VSS.n4255 VSS.n4254 0.0405
R23521 VSS.n3463 VSS.n3462 0.0405
R23522 VSS.n3462 VSS.n3461 0.0405
R23523 VSS.n3461 VSS.n3200 0.0405
R23524 VSS.n3457 VSS.n3200 0.0405
R23525 VSS.n3457 VSS.n3456 0.0405
R23526 VSS.n3456 VSS.n3455 0.0405
R23527 VSS.n3455 VSS.n3205 0.0405
R23528 VSS.n3451 VSS.n3205 0.0405
R23529 VSS.n3451 VSS.n3450 0.0405
R23530 VSS.n3450 VSS.n3449 0.0405
R23531 VSS.n3449 VSS.n3445 0.0405
R23532 VSS.n3445 VSS.n2926 0.0405
R23533 VSS.n3695 VSS.n3079 0.0405
R23534 VSS.n3720 VSS.n3079 0.0405
R23535 VSS.n3720 VSS.n3076 0.0405
R23536 VSS.n3725 VSS.n3076 0.0405
R23537 VSS.n3725 VSS.n3077 0.0405
R23538 VSS.n3077 VSS.n3065 0.0405
R23539 VSS.n3753 VSS.n3065 0.0405
R23540 VSS.n3753 VSS.n3062 0.0405
R23541 VSS.n3758 VSS.n3062 0.0405
R23542 VSS.n3758 VSS.n3063 0.0405
R23543 VSS.n3063 VSS.n3046 0.0405
R23544 VSS.n3777 VSS.n3046 0.0405
R23545 VSS.n3777 VSS.n3044 0.0405
R23546 VSS.n3781 VSS.n3044 0.0405
R23547 VSS.n3801 VSS.n3037 0.0405
R23548 VSS.n3801 VSS.n3034 0.0405
R23549 VSS.n3808 VSS.n3034 0.0405
R23550 VSS.n3808 VSS.n3035 0.0405
R23551 VSS.n3804 VSS.n3035 0.0405
R23552 VSS.n3804 VSS.n3020 0.0405
R23553 VSS.n3839 VSS.n3020 0.0405
R23554 VSS.n3839 VSS.n3018 0.0405
R23555 VSS.n3843 VSS.n3018 0.0405
R23556 VSS.n3843 VSS.n3008 0.0405
R23557 VSS.n4196 VSS.n3008 0.0405
R23558 VSS.n4196 VSS.n3005 0.0405
R23559 VSS.n3694 VSS.n3078 0.0405
R23560 VSS.n3721 VSS.n3078 0.0405
R23561 VSS.n3722 VSS.n3721 0.0405
R23562 VSS.n3724 VSS.n3722 0.0405
R23563 VSS.n3724 VSS.n3723 0.0405
R23564 VSS.n3723 VSS.n3064 0.0405
R23565 VSS.n3754 VSS.n3064 0.0405
R23566 VSS.n3755 VSS.n3754 0.0405
R23567 VSS.n3757 VSS.n3755 0.0405
R23568 VSS.n3757 VSS.n3756 0.0405
R23569 VSS.n3756 VSS.n3045 0.0405
R23570 VSS.n3778 VSS.n3045 0.0405
R23571 VSS.n3779 VSS.n3778 0.0405
R23572 VSS.n3780 VSS.n3779 0.0405
R23573 VSS.n3802 VSS.n3036 0.0405
R23574 VSS.n3803 VSS.n3802 0.0405
R23575 VSS.n3807 VSS.n3803 0.0405
R23576 VSS.n3807 VSS.n3806 0.0405
R23577 VSS.n3806 VSS.n3805 0.0405
R23578 VSS.n3805 VSS.n3019 0.0405
R23579 VSS.n3840 VSS.n3019 0.0405
R23580 VSS.n3841 VSS.n3840 0.0405
R23581 VSS.n3842 VSS.n3841 0.0405
R23582 VSS.n3842 VSS.n3007 0.0405
R23583 VSS.n4197 VSS.n3007 0.0405
R23584 VSS.n4198 VSS.n4197 0.0405
R23585 VSS.n3464 VSS.n3196 0.0405
R23586 VSS.n3460 VSS.n3196 0.0405
R23587 VSS.n3460 VSS.n3459 0.0405
R23588 VSS.n3459 VSS.n3458 0.0405
R23589 VSS.n3458 VSS.n3201 0.0405
R23590 VSS.n3454 VSS.n3201 0.0405
R23591 VSS.n3454 VSS.n3453 0.0405
R23592 VSS.n3453 VSS.n3452 0.0405
R23593 VSS.n3452 VSS.n3206 0.0405
R23594 VSS.n3448 VSS.n3206 0.0405
R23595 VSS.n3448 VSS.n3447 0.0405
R23596 VSS.n3447 VSS.n3446 0.0405
R23597 VSS.n2951 VSS.n2950 0.0405
R23598 VSS.n4265 VSS.n2951 0.0405
R23599 VSS.n4265 VSS.n4264 0.0405
R23600 VSS.n4264 VSS.n4263 0.0405
R23601 VSS.n4263 VSS.n2952 0.0405
R23602 VSS.n4259 VSS.n2952 0.0405
R23603 VSS.n4259 VSS.n4258 0.0405
R23604 VSS.n4258 VSS.n4257 0.0405
R23605 VSS.n4257 VSS.n2957 0.0405
R23606 VSS.n4253 VSS.n2957 0.0405
R23607 VSS.n2739 VSS.n2738 0.0405
R23608 VSS.n2738 VSS.n2737 0.0405
R23609 VSS.n2737 VSS.n1493 0.0405
R23610 VSS.n2733 VSS.n1493 0.0405
R23611 VSS.n2733 VSS.n2732 0.0405
R23612 VSS.n2732 VSS.n2731 0.0405
R23613 VSS.n2731 VSS.n1498 0.0405
R23614 VSS.n2727 VSS.n1498 0.0405
R23615 VSS.n2727 VSS.n2726 0.0405
R23616 VSS.n2726 VSS.n2725 0.0405
R23617 VSS.n2725 VSS.n1503 0.0405
R23618 VSS.n2721 VSS.n1503 0.0405
R23619 VSS.n2721 VSS.n2720 0.0405
R23620 VSS.n2720 VSS.n2719 0.0405
R23621 VSS.n2715 VSS.n1508 0.0405
R23622 VSS.n2715 VSS.n2714 0.0405
R23623 VSS.n2714 VSS.n2713 0.0405
R23624 VSS.n2713 VSS.n1513 0.0405
R23625 VSS.n2709 VSS.n1513 0.0405
R23626 VSS.n2709 VSS.n2708 0.0405
R23627 VSS.n2708 VSS.n2707 0.0405
R23628 VSS.n2707 VSS.n1518 0.0405
R23629 VSS.n2703 VSS.n1518 0.0405
R23630 VSS.n2703 VSS.n2702 0.0405
R23631 VSS.n2702 VSS.n2701 0.0405
R23632 VSS.n2701 VSS.n1523 0.0405
R23633 VSS.n2740 VSS.n1489 0.0405
R23634 VSS.n2736 VSS.n1489 0.0405
R23635 VSS.n2736 VSS.n2735 0.0405
R23636 VSS.n2735 VSS.n2734 0.0405
R23637 VSS.n2734 VSS.n1494 0.0405
R23638 VSS.n2730 VSS.n1494 0.0405
R23639 VSS.n2730 VSS.n2729 0.0405
R23640 VSS.n2729 VSS.n2728 0.0405
R23641 VSS.n2728 VSS.n1499 0.0405
R23642 VSS.n2724 VSS.n1499 0.0405
R23643 VSS.n2724 VSS.n2723 0.0405
R23644 VSS.n2723 VSS.n2722 0.0405
R23645 VSS.n2722 VSS.n1504 0.0405
R23646 VSS.n2718 VSS.n1504 0.0405
R23647 VSS.n2717 VSS.n2716 0.0405
R23648 VSS.n2716 VSS.n1509 0.0405
R23649 VSS.n2712 VSS.n1509 0.0405
R23650 VSS.n2712 VSS.n2711 0.0405
R23651 VSS.n2711 VSS.n2710 0.0405
R23652 VSS.n2710 VSS.n1514 0.0405
R23653 VSS.n2706 VSS.n1514 0.0405
R23654 VSS.n2706 VSS.n2705 0.0405
R23655 VSS.n2705 VSS.n2704 0.0405
R23656 VSS.n2704 VSS.n1519 0.0405
R23657 VSS.n2700 VSS.n1519 0.0405
R23658 VSS.n2700 VSS.n2699 0.0405
R23659 VSS.n2186 VSS.n2026 0.0405
R23660 VSS.n2186 VSS.n2027 0.0405
R23661 VSS.n2182 VSS.n2027 0.0405
R23662 VSS.n2182 VSS.n2181 0.0405
R23663 VSS.n2181 VSS.n2180 0.0405
R23664 VSS.n2180 VSS.n2177 0.0405
R23665 VSS.n2177 VSS.n1984 0.0405
R23666 VSS.n2279 VSS.n1984 0.0405
R23667 VSS.n2279 VSS.n1979 0.0405
R23668 VSS.n2284 VSS.n1979 0.0405
R23669 VSS.n2284 VSS.n1982 0.0405
R23670 VSS.n1982 VSS.n1959 0.0405
R23671 VSS.n2332 VSS.n1959 0.0405
R23672 VSS.n2332 VSS.n1957 0.0405
R23673 VSS.n2336 VSS.n1940 0.0405
R23674 VSS.n2375 VSS.n1940 0.0405
R23675 VSS.n2375 VSS.n1937 0.0405
R23676 VSS.n2384 VSS.n1937 0.0405
R23677 VSS.n2384 VSS.n1938 0.0405
R23678 VSS.n2380 VSS.n1938 0.0405
R23679 VSS.n2380 VSS.n2379 0.0405
R23680 VSS.n2379 VSS.n1906 0.0405
R23681 VSS.n2467 VSS.n1906 0.0405
R23682 VSS.n2467 VSS.n1904 0.0405
R23683 VSS.n2471 VSS.n1904 0.0405
R23684 VSS.n2471 VSS.n1892 0.0405
R23685 VSS.n2185 VSS.n2175 0.0405
R23686 VSS.n2185 VSS.n2184 0.0405
R23687 VSS.n2184 VSS.n2183 0.0405
R23688 VSS.n2183 VSS.n2176 0.0405
R23689 VSS.n2179 VSS.n2176 0.0405
R23690 VSS.n2179 VSS.n2178 0.0405
R23691 VSS.n2178 VSS.n1983 0.0405
R23692 VSS.n2280 VSS.n1983 0.0405
R23693 VSS.n2281 VSS.n2280 0.0405
R23694 VSS.n2283 VSS.n2281 0.0405
R23695 VSS.n2283 VSS.n2282 0.0405
R23696 VSS.n2282 VSS.n1958 0.0405
R23697 VSS.n2333 VSS.n1958 0.0405
R23698 VSS.n2334 VSS.n2333 0.0405
R23699 VSS.n2335 VSS.n1939 0.0405
R23700 VSS.n2376 VSS.n1939 0.0405
R23701 VSS.n2377 VSS.n2376 0.0405
R23702 VSS.n2383 VSS.n2377 0.0405
R23703 VSS.n2383 VSS.n2382 0.0405
R23704 VSS.n2382 VSS.n2381 0.0405
R23705 VSS.n2381 VSS.n2378 0.0405
R23706 VSS.n2378 VSS.n1905 0.0405
R23707 VSS.n2468 VSS.n1905 0.0405
R23708 VSS.n2469 VSS.n2468 0.0405
R23709 VSS.n2470 VSS.n2469 0.0405
R23710 VSS.n2470 VSS.n1891 0.0405
R23711 VSS.n1088 VSS.n449 0.0403551
R23712 VSS.n1421 VSS.n127 0.0400614
R23713 VSS.n242 VSS.n142 0.0400614
R23714 VSS.n262 VSS.n133 0.0400614
R23715 VSS.n1371 VSS.n331 0.0400614
R23716 VSS.n1357 VSS.n312 0.0400614
R23717 VSS.n1331 VSS.n1330 0.0400614
R23718 VSS.n2900 VSS.n39 0.039
R23719 VSS.n864 VSS.n863 0.0384472
R23720 VSS.n880 VSS.n879 0.0384472
R23721 VSS.n1213 VSS.n1212 0.0384472
R23722 VSS.n415 VSS.n414 0.0384472
R23723 VSS.n240 VSS.n129 0.0381316
R23724 VSS.n264 VSS.n137 0.0381316
R23725 VSS.n1373 VSS.n308 0.0381316
R23726 VSS.n1355 VSS.n324 0.0381316
R23727 VSS.n1214 VSS 0.038
R23728 VSS VSS.n1180 0.038
R23729 VSS VSS.n413 0.038
R23730 VSS.n1250 VSS 0.038
R23731 VSS.n238 VSS.n153 0.0362018
R23732 VSS.n170 VSS.n134 0.0362018
R23733 VSS.n1377 VSS.n1376 0.0362018
R23734 VSS.n1353 VSS.n313 0.0362018
R23735 VSS.n3781 VSS.n3037 0.0360676
R23736 VSS.n3780 VSS.n3036 0.0360676
R23737 VSS.n3467 VSS.n3466 0.0360676
R23738 VSS.n3467 VSS.n3183 0.0360676
R23739 VSS.n3492 VSS.n3183 0.0360676
R23740 VSS.n3493 VSS.n3492 0.0360676
R23741 VSS.n3494 VSS.n3493 0.0360676
R23742 VSS.n3494 VSS.n3170 0.0360676
R23743 VSS.n3517 VSS.n3170 0.0360676
R23744 VSS.n3518 VSS.n3517 0.0360676
R23745 VSS.n3519 VSS.n3518 0.0360676
R23746 VSS.n3520 VSS.n3519 0.0360676
R23747 VSS.n3521 VSS.n3520 0.0360676
R23748 VSS.n3521 VSS.n3151 0.0360676
R23749 VSS.n3563 VSS.n3151 0.0360676
R23750 VSS.n3564 VSS.n3563 0.0360676
R23751 VSS.n3565 VSS.n3564 0.0360676
R23752 VSS.n3565 VSS.n3134 0.0360676
R23753 VSS.n3583 VSS.n3134 0.0360676
R23754 VSS.n3584 VSS.n3583 0.0360676
R23755 VSS.n3585 VSS.n3584 0.0360676
R23756 VSS.n3586 VSS.n3585 0.0360676
R23757 VSS.n3587 VSS.n3586 0.0360676
R23758 VSS.n3587 VSS.n3116 0.0360676
R23759 VSS.n3624 VSS.n3116 0.0360676
R23760 VSS.n3625 VSS.n3624 0.0360676
R23761 VSS.n3626 VSS.n3625 0.0360676
R23762 VSS.n3627 VSS.n3626 0.0360676
R23763 VSS.n3628 VSS.n3627 0.0360676
R23764 VSS.n3628 VSS.n3099 0.0360676
R23765 VSS.n3673 VSS.n3099 0.0360676
R23766 VSS.n3674 VSS.n3673 0.0360676
R23767 VSS.n3675 VSS.n3674 0.0360676
R23768 VSS.n3675 VSS.n3090 0.0360676
R23769 VSS.n3692 VSS.n3090 0.0360676
R23770 VSS.n3469 VSS.n3468 0.0360676
R23771 VSS.n3468 VSS.n3184 0.0360676
R23772 VSS.n3491 VSS.n3184 0.0360676
R23773 VSS.n3491 VSS.n3182 0.0360676
R23774 VSS.n3495 VSS.n3182 0.0360676
R23775 VSS.n3495 VSS.n3171 0.0360676
R23776 VSS.n3516 VSS.n3171 0.0360676
R23777 VSS.n3516 VSS.n3169 0.0360676
R23778 VSS.n3530 VSS.n3169 0.0360676
R23779 VSS.n3530 VSS.n3529 0.0360676
R23780 VSS.n3529 VSS.n3522 0.0360676
R23781 VSS.n3522 VSS.n3152 0.0360676
R23782 VSS.n3562 VSS.n3152 0.0360676
R23783 VSS.n3562 VSS.n3150 0.0360676
R23784 VSS.n3566 VSS.n3150 0.0360676
R23785 VSS.n3566 VSS.n3135 0.0360676
R23786 VSS.n3582 VSS.n3135 0.0360676
R23787 VSS.n3582 VSS.n3133 0.0360676
R23788 VSS.n3596 VSS.n3133 0.0360676
R23789 VSS.n3596 VSS.n3595 0.0360676
R23790 VSS.n3595 VSS.n3588 0.0360676
R23791 VSS.n3588 VSS.n3117 0.0360676
R23792 VSS.n3623 VSS.n3117 0.0360676
R23793 VSS.n3623 VSS.n3115 0.0360676
R23794 VSS.n3631 VSS.n3115 0.0360676
R23795 VSS.n3631 VSS.n3630 0.0360676
R23796 VSS.n3630 VSS.n3629 0.0360676
R23797 VSS.n3629 VSS.n3100 0.0360676
R23798 VSS.n3672 VSS.n3100 0.0360676
R23799 VSS.n3672 VSS.n3098 0.0360676
R23800 VSS.n3676 VSS.n3098 0.0360676
R23801 VSS.n3676 VSS.n3091 0.0360676
R23802 VSS.n3691 VSS.n3091 0.0360676
R23803 VSS.n4250 VSS.n4249 0.0360676
R23804 VSS.n4249 VSS.n4248 0.0360676
R23805 VSS.n4248 VSS.n2966 0.0360676
R23806 VSS.n4244 VSS.n2966 0.0360676
R23807 VSS.n4244 VSS.n4243 0.0360676
R23808 VSS.n4243 VSS.n4242 0.0360676
R23809 VSS.n4242 VSS.n2971 0.0360676
R23810 VSS.n4238 VSS.n2971 0.0360676
R23811 VSS.n4238 VSS.n4237 0.0360676
R23812 VSS.n4237 VSS.n4236 0.0360676
R23813 VSS.n4236 VSS.n2976 0.0360676
R23814 VSS.n4232 VSS.n2976 0.0360676
R23815 VSS.n4232 VSS.n4231 0.0360676
R23816 VSS.n4231 VSS.n4230 0.0360676
R23817 VSS.n4230 VSS.n2981 0.0360676
R23818 VSS.n4226 VSS.n2981 0.0360676
R23819 VSS.n4226 VSS.n4225 0.0360676
R23820 VSS.n4225 VSS.n4224 0.0360676
R23821 VSS.n4224 VSS.n2986 0.0360676
R23822 VSS.n4220 VSS.n2986 0.0360676
R23823 VSS.n4220 VSS.n4219 0.0360676
R23824 VSS.n4219 VSS.n4218 0.0360676
R23825 VSS.n4218 VSS.n2991 0.0360676
R23826 VSS.n4214 VSS.n2991 0.0360676
R23827 VSS.n4214 VSS.n4213 0.0360676
R23828 VSS.n4213 VSS.n4212 0.0360676
R23829 VSS.n4212 VSS.n2996 0.0360676
R23830 VSS.n4208 VSS.n2996 0.0360676
R23831 VSS.n4208 VSS.n4207 0.0360676
R23832 VSS.n4207 VSS.n4206 0.0360676
R23833 VSS.n4206 VSS.n3001 0.0360676
R23834 VSS.n4202 VSS.n3001 0.0360676
R23835 VSS.n4202 VSS.n4201 0.0360676
R23836 VSS.n4251 VSS.n2962 0.0360676
R23837 VSS.n4247 VSS.n2962 0.0360676
R23838 VSS.n4247 VSS.n4246 0.0360676
R23839 VSS.n4246 VSS.n4245 0.0360676
R23840 VSS.n4245 VSS.n2967 0.0360676
R23841 VSS.n4241 VSS.n2967 0.0360676
R23842 VSS.n4241 VSS.n4240 0.0360676
R23843 VSS.n4240 VSS.n4239 0.0360676
R23844 VSS.n4239 VSS.n2972 0.0360676
R23845 VSS.n4235 VSS.n2972 0.0360676
R23846 VSS.n4235 VSS.n4234 0.0360676
R23847 VSS.n4234 VSS.n4233 0.0360676
R23848 VSS.n4233 VSS.n2977 0.0360676
R23849 VSS.n4229 VSS.n2977 0.0360676
R23850 VSS.n4229 VSS.n4228 0.0360676
R23851 VSS.n4228 VSS.n4227 0.0360676
R23852 VSS.n4227 VSS.n2982 0.0360676
R23853 VSS.n4223 VSS.n2982 0.0360676
R23854 VSS.n4223 VSS.n4222 0.0360676
R23855 VSS.n4222 VSS.n4221 0.0360676
R23856 VSS.n4221 VSS.n2987 0.0360676
R23857 VSS.n4217 VSS.n2987 0.0360676
R23858 VSS.n4217 VSS.n4216 0.0360676
R23859 VSS.n4216 VSS.n4215 0.0360676
R23860 VSS.n4215 VSS.n2992 0.0360676
R23861 VSS.n4211 VSS.n2992 0.0360676
R23862 VSS.n4211 VSS.n4210 0.0360676
R23863 VSS.n4210 VSS.n4209 0.0360676
R23864 VSS.n4209 VSS.n2997 0.0360676
R23865 VSS.n4205 VSS.n2997 0.0360676
R23866 VSS.n4205 VSS.n4204 0.0360676
R23867 VSS.n4204 VSS.n4203 0.0360676
R23868 VSS.n4203 VSS.n3002 0.0360676
R23869 VSS.n2719 VSS.n1508 0.0360676
R23870 VSS.n2718 VSS.n2717 0.0360676
R23871 VSS.n2336 VSS.n1957 0.0360676
R23872 VSS.n2335 VSS.n2334 0.0360676
R23873 VSS.n2508 VSS.n2507 0.0360676
R23874 VSS.n2508 VSS.n1881 0.0360676
R23875 VSS.n2528 VSS.n1881 0.0360676
R23876 VSS.n2529 VSS.n2528 0.0360676
R23877 VSS.n2530 VSS.n2529 0.0360676
R23878 VSS.n2530 VSS.n1867 0.0360676
R23879 VSS.n2551 VSS.n1867 0.0360676
R23880 VSS.n2552 VSS.n2551 0.0360676
R23881 VSS.n2553 VSS.n2552 0.0360676
R23882 VSS.n2554 VSS.n2553 0.0360676
R23883 VSS.n2554 VSS.n1855 0.0360676
R23884 VSS.n2582 VSS.n1855 0.0360676
R23885 VSS.n2583 VSS.n2582 0.0360676
R23886 VSS.n2584 VSS.n2583 0.0360676
R23887 VSS.n2585 VSS.n2584 0.0360676
R23888 VSS.n2585 VSS.n1838 0.0360676
R23889 VSS.n2606 VSS.n1838 0.0360676
R23890 VSS.n2607 VSS.n2606 0.0360676
R23891 VSS.n2608 VSS.n2607 0.0360676
R23892 VSS.n2608 VSS.n1828 0.0360676
R23893 VSS.n2629 VSS.n1828 0.0360676
R23894 VSS.n2630 VSS.n2629 0.0360676
R23895 VSS.n2631 VSS.n2630 0.0360676
R23896 VSS.n2632 VSS.n2631 0.0360676
R23897 VSS.n2632 VSS.n1817 0.0360676
R23898 VSS.n2660 VSS.n1817 0.0360676
R23899 VSS.n2661 VSS.n2660 0.0360676
R23900 VSS.n2662 VSS.n2661 0.0360676
R23901 VSS.n2662 VSS.n1808 0.0360676
R23902 VSS.n2684 VSS.n1808 0.0360676
R23903 VSS.n2685 VSS.n2684 0.0360676
R23904 VSS.n2686 VSS.n2685 0.0360676
R23905 VSS.n2686 VSS.n1524 0.0360676
R23906 VSS.n2509 VSS.n1890 0.0360676
R23907 VSS.n2509 VSS.n1882 0.0360676
R23908 VSS.n2527 VSS.n1882 0.0360676
R23909 VSS.n2527 VSS.n1880 0.0360676
R23910 VSS.n2531 VSS.n1880 0.0360676
R23911 VSS.n2531 VSS.n1868 0.0360676
R23912 VSS.n2550 VSS.n1868 0.0360676
R23913 VSS.n2550 VSS.n1866 0.0360676
R23914 VSS.n2556 VSS.n1866 0.0360676
R23915 VSS.n2556 VSS.n2555 0.0360676
R23916 VSS.n2555 VSS.n1856 0.0360676
R23917 VSS.n2581 VSS.n1856 0.0360676
R23918 VSS.n2581 VSS.n1854 0.0360676
R23919 VSS.n2587 VSS.n1854 0.0360676
R23920 VSS.n2587 VSS.n2586 0.0360676
R23921 VSS.n2586 VSS.n1839 0.0360676
R23922 VSS.n2605 VSS.n1839 0.0360676
R23923 VSS.n2605 VSS.n1837 0.0360676
R23924 VSS.n2609 VSS.n1837 0.0360676
R23925 VSS.n2609 VSS.n1829 0.0360676
R23926 VSS.n2628 VSS.n1829 0.0360676
R23927 VSS.n2628 VSS.n1827 0.0360676
R23928 VSS.n2634 VSS.n1827 0.0360676
R23929 VSS.n2634 VSS.n2633 0.0360676
R23930 VSS.n2633 VSS.n1818 0.0360676
R23931 VSS.n2659 VSS.n1818 0.0360676
R23932 VSS.n2659 VSS.n1816 0.0360676
R23933 VSS.n2663 VSS.n1816 0.0360676
R23934 VSS.n2663 VSS.n1809 0.0360676
R23935 VSS.n2683 VSS.n1809 0.0360676
R23936 VSS.n2683 VSS.n1807 0.0360676
R23937 VSS.n2687 VSS.n1807 0.0360676
R23938 VSS.n2687 VSS.n1525 0.0360676
R23939 VSS.n2161 VSS.n2029 0.0360676
R23940 VSS.n2161 VSS.n2057 0.0360676
R23941 VSS.n2157 VSS.n2057 0.0360676
R23942 VSS.n2157 VSS.n2156 0.0360676
R23943 VSS.n2156 VSS.n2155 0.0360676
R23944 VSS.n2155 VSS.n2062 0.0360676
R23945 VSS.n2151 VSS.n2062 0.0360676
R23946 VSS.n2151 VSS.n2150 0.0360676
R23947 VSS.n2150 VSS.n2149 0.0360676
R23948 VSS.n2149 VSS.n2067 0.0360676
R23949 VSS.n2145 VSS.n2067 0.0360676
R23950 VSS.n2145 VSS.n1441 0.0360676
R23951 VSS.n1470 VSS.n1442 0.0360676
R23952 VSS.n2761 VSS.n1470 0.0360676
R23953 VSS.n2761 VSS.n1471 0.0360676
R23954 VSS.n2757 VSS.n1471 0.0360676
R23955 VSS.n2757 VSS.n2756 0.0360676
R23956 VSS.n2756 VSS.n2755 0.0360676
R23957 VSS.n2755 VSS.n1478 0.0360676
R23958 VSS.n2751 VSS.n1478 0.0360676
R23959 VSS.n2751 VSS.n2750 0.0360676
R23960 VSS.n2750 VSS.n2749 0.0360676
R23961 VSS.n2749 VSS.n1483 0.0360676
R23962 VSS.n2745 VSS.n1483 0.0360676
R23963 VSS.n2745 VSS.n2744 0.0360676
R23964 VSS.n2744 VSS.n2743 0.0360676
R23965 VSS.n2160 VSS.n2028 0.0360676
R23966 VSS.n2160 VSS.n2159 0.0360676
R23967 VSS.n2159 VSS.n2158 0.0360676
R23968 VSS.n2158 VSS.n2058 0.0360676
R23969 VSS.n2154 VSS.n2058 0.0360676
R23970 VSS.n2154 VSS.n2153 0.0360676
R23971 VSS.n2153 VSS.n2152 0.0360676
R23972 VSS.n2152 VSS.n2063 0.0360676
R23973 VSS.n2148 VSS.n2063 0.0360676
R23974 VSS.n2148 VSS.n2147 0.0360676
R23975 VSS.n2147 VSS.n2146 0.0360676
R23976 VSS.n2146 VSS.n2068 0.0360676
R23977 VSS.n1473 VSS.n1472 0.0360676
R23978 VSS.n2760 VSS.n1473 0.0360676
R23979 VSS.n2760 VSS.n2759 0.0360676
R23980 VSS.n2759 VSS.n2758 0.0360676
R23981 VSS.n2758 VSS.n1474 0.0360676
R23982 VSS.n2754 VSS.n1474 0.0360676
R23983 VSS.n2754 VSS.n2753 0.0360676
R23984 VSS.n2753 VSS.n2752 0.0360676
R23985 VSS.n2752 VSS.n1479 0.0360676
R23986 VSS.n2748 VSS.n1479 0.0360676
R23987 VSS.n2748 VSS.n2747 0.0360676
R23988 VSS.n2747 VSS.n2746 0.0360676
R23989 VSS.n2746 VSS.n1484 0.0360676
R23990 VSS.n2742 VSS.n1484 0.0360676
R23991 VSS.n1147 VSS.n1146 0.0351579
R23992 VSS.n1152 VSS.n1151 0.0351579
R23993 VSS.n185 VSS.n152 0.0342719
R23994 VSS.n272 VSS.n136 0.0342719
R23995 VSS.n1416 VSS.n158 0.0342719
R23996 VSS.n1379 VSS.n307 0.0342719
R23997 VSS.n1351 VSS.n323 0.0342719
R23998 VSS.n1440 VSS.n109 0.0342165
R23999 VSS.n198 VSS.n109 0.0342165
R24000 VSS.n199 VSS.n198 0.0342165
R24001 VSS.n200 VSS.n199 0.0342165
R24002 VSS.n202 VSS.n200 0.0342165
R24003 VSS.n203 VSS.n202 0.0342165
R24004 VSS.n204 VSS.n203 0.0342165
R24005 VSS.n205 VSS.n204 0.0342165
R24006 VSS.n207 VSS.n205 0.0342165
R24007 VSS.n208 VSS.n207 0.0342165
R24008 VSS.n209 VSS.n208 0.0342165
R24009 VSS.n210 VSS.n209 0.0342165
R24010 VSS.n212 VSS.n210 0.0342165
R24011 VSS.n213 VSS.n212 0.0342165
R24012 VSS.n214 VSS.n213 0.0342165
R24013 VSS.n214 VSS.n193 0.0342165
R24014 VSS.n223 VSS.n193 0.0342165
R24015 VSS.n224 VSS.n223 0.0342165
R24016 VSS.n225 VSS.n224 0.0342165
R24017 VSS.n225 VSS.n188 0.0342165
R24018 VSS.n234 VSS.n188 0.0342165
R24019 VSS.n235 VSS.n234 0.0342165
R24020 VSS.n236 VSS.n235 0.0342165
R24021 VSS.n236 VSS.n183 0.0342165
R24022 VSS.n245 VSS.n183 0.0342165
R24023 VSS.n246 VSS.n245 0.0342165
R24024 VSS.n247 VSS.n246 0.0342165
R24025 VSS.n247 VSS.n178 0.0342165
R24026 VSS.n256 VSS.n178 0.0342165
R24027 VSS.n257 VSS.n256 0.0342165
R24028 VSS.n258 VSS.n257 0.0342165
R24029 VSS.n258 VSS.n173 0.0342165
R24030 VSS.n267 VSS.n173 0.0342165
R24031 VSS.n268 VSS.n267 0.0342165
R24032 VSS.n270 VSS.n268 0.0342165
R24033 VSS.n270 VSS.n269 0.0342165
R24034 VSS.n269 VSS.n168 0.0342165
R24035 VSS.n280 VSS.n168 0.0342165
R24036 VSS.n281 VSS.n280 0.0342165
R24037 VSS.n282 VSS.n281 0.0342165
R24038 VSS.n283 VSS.n282 0.0342165
R24039 VSS.n285 VSS.n283 0.0342165
R24040 VSS.n286 VSS.n285 0.0342165
R24041 VSS.n287 VSS.n286 0.0342165
R24042 VSS.n288 VSS.n287 0.0342165
R24043 VSS.n1400 VSS.n288 0.0342165
R24044 VSS.n1399 VSS.n289 0.0342165
R24045 VSS.n1264 VSS.n289 0.0342165
R24046 VSS.n1265 VSS.n1264 0.0342165
R24047 VSS.n1267 VSS.n1265 0.0342165
R24048 VSS.n1268 VSS.n1267 0.0342165
R24049 VSS.n1269 VSS.n1268 0.0342165
R24050 VSS.n1271 VSS.n1269 0.0342165
R24051 VSS.n1272 VSS.n1271 0.0342165
R24052 VSS.n1273 VSS.n1272 0.0342165
R24053 VSS.n1274 VSS.n1273 0.0342165
R24054 VSS.n1276 VSS.n1274 0.0342165
R24055 VSS.n1277 VSS.n1276 0.0342165
R24056 VSS.n1278 VSS.n1277 0.0342165
R24057 VSS.n1279 VSS.n1278 0.0342165
R24058 VSS.n1280 VSS.n1279 0.0342165
R24059 VSS.n1281 VSS.n1280 0.0342165
R24060 VSS.n1282 VSS.n1281 0.0342165
R24061 VSS.n1283 VSS.n1282 0.0342165
R24062 VSS.n1284 VSS.n1283 0.0342165
R24063 VSS.n1285 VSS.n1284 0.0342165
R24064 VSS.n1286 VSS.n1285 0.0342165
R24065 VSS.n1287 VSS.n1286 0.0342165
R24066 VSS.n1288 VSS.n1287 0.0342165
R24067 VSS.n1289 VSS.n1288 0.0342165
R24068 VSS.n1290 VSS.n1289 0.0342165
R24069 VSS.n1291 VSS.n1290 0.0342165
R24070 VSS.n1292 VSS.n1291 0.0342165
R24071 VSS.n1293 VSS.n1292 0.0342165
R24072 VSS.n1294 VSS.n1293 0.0342165
R24073 VSS.n1295 VSS.n1294 0.0342165
R24074 VSS.n1296 VSS.n1295 0.0342165
R24075 VSS.n1297 VSS.n1296 0.0342165
R24076 VSS.n1298 VSS.n1297 0.0342165
R24077 VSS.n1299 VSS.n1298 0.0342165
R24078 VSS.n1319 VSS.n1300 0.0342165
R24079 VSS.n1319 VSS.n1318 0.0342165
R24080 VSS.n1318 VSS.n1317 0.0342165
R24081 VSS.n1317 VSS.n1301 0.0342165
R24082 VSS.n1313 VSS.n1301 0.0342165
R24083 VSS.n708 VSS.n707 0.0333479
R24084 VSS.n713 VSS.n708 0.0326581
R24085 VSS.n734 VSS.n733 0.0324848
R24086 VSS.n1421 VSS.n1420 0.0323421
R24087 VSS.n231 VSS.n151 0.0323421
R24088 VSS.n274 VSS.n135 0.0323421
R24089 VSS.n1415 VSS.n156 0.0323421
R24090 VSS.n1387 VSS.n300 0.0323421
R24091 VSS.n1380 VSS.n306 0.0323421
R24092 VSS.n1349 VSS.n314 0.0323421
R24093 VSS.n962 VSS.n516 0.0319824
R24094 VSS.n796 VSS.n787 0.031863
R24095 VSS.n878 VSS.n877 0.031863
R24096 VSS.n2895 VSS.n46 0.0316667
R24097 VSS.n835 VSS.n834 0.0309472
R24098 VSS.n786 VSS.n785 0.0309472
R24099 VSS.n833 VSS.n832 0.0309472
R24100 VSS.n923 VSS.n922 0.0309472
R24101 VSS.n782 VSS.n781 0.0309472
R24102 VSS.n913 VSS.n912 0.0309472
R24103 VSS.n1189 VSS.n1188 0.0309472
R24104 VSS.n1182 VSS.n1181 0.0309472
R24105 VSS.n1242 VSS.n1241 0.0309472
R24106 VSS.n1249 VSS.n1248 0.0309472
R24107 VSS.n833 VSS 0.0305
R24108 VSS VSS.n862 0.0305
R24109 VSS.n785 VSS 0.0305
R24110 VSS.n912 VSS 0.0305
R24111 VSS.n896 VSS 0.0305
R24112 VSS.n782 VSS 0.0305
R24113 VSS.n1181 VSS 0.0305
R24114 VSS VSS.n1249 0.0305
R24115 VSS.n144 VSS.n128 0.0304123
R24116 VSS.n229 VSS.n150 0.0304123
R24117 VSS.n1412 VSS.n157 0.0304123
R24118 VSS.n1388 VSS.n296 0.0304123
R24119 VSS.n1347 VSS.n322 0.0304123
R24120 VSS.n1333 VSS.n319 0.0304123
R24121 VSS.n2888 VSS.n32 0.0298333
R24122 VSS.n1256 VSS 0.0291391
R24123 VSS.n195 VSS.n145 0.0284825
R24124 VSS.n227 VSS.n149 0.0284825
R24125 VSS.n1345 VSS.n315 0.0284825
R24126 VSS.n1335 VSS.n317 0.0284825
R24127 VSS.n748 VSS 0.028469
R24128 VSS.n1257 VSS.n356 0.0281035
R24129 VSS.n2844 VSS.n2843 0.028
R24130 VSS.n843 VSS.n842 0.0266282
R24131 VSS.n1250 VSS.n362 0.0266282
R24132 VSS.n216 VSS.n146 0.0265526
R24133 VSS.n190 VSS.n148 0.0265526
R24134 VSS.n1343 VSS.n321 0.0265526
R24135 VSS.n1337 VSS.n320 0.0265526
R24136 VSS.n357 VSS.n356 0.0261075
R24137 VSS.n251 VSS.n140 0.0250913
R24138 VSS.n253 VSS.n140 0.0250913
R24139 VSS.n1365 VSS.n329 0.0250913
R24140 VSS.n1363 VSS.n329 0.0250913
R24141 VSS.n746 VSS.n745 0.0249824
R24142 VSS.n218 VSS.n147 0.0246228
R24143 VSS.n220 VSS.n147 0.0246228
R24144 VSS.n1341 VSS.n316 0.0246228
R24145 VSS.n1339 VSS.n316 0.0246228
R24146 VSS.n1385 VSS 0.0236579
R24147 VSS VSS.n318 0.0236579
R24148 VSS.n3463 VSS.n3195 0.0234189
R24149 VSS.n3695 VSS.n3089 0.0234189
R24150 VSS.n3694 VSS.n3693 0.0234189
R24151 VSS.n3465 VSS.n3464 0.0234189
R24152 VSS.n2739 VSS.n1488 0.0234189
R24153 VSS.n2741 VSS.n2740 0.0234189
R24154 VSS.n2173 VSS.n2026 0.0234189
R24155 VSS.n2175 VSS.n2174 0.0234189
R24156 VSS.n4254 VSS.n2961 0.0233108
R24157 VSS.n4200 VSS.n3005 0.0233108
R24158 VSS.n4199 VSS.n4198 0.0233108
R24159 VSS.n4253 VSS.n4252 0.0233108
R24160 VSS.n2697 VSS.n1523 0.0233108
R24161 VSS.n2699 VSS.n2698 0.0233108
R24162 VSS.n2505 VSS.n1892 0.0233108
R24163 VSS.n2506 VSS.n1891 0.0233108
R24164 VSS VSS.n864 0.023
R24165 VSS.n879 VSS 0.023
R24166 VSS VSS.n1213 0.023
R24167 VSS.n1191 VSS 0.023
R24168 VSS.n414 VSS 0.023
R24169 VSS VSS.n1239 0.023
R24170 VSS.n3466 VSS.n3465 0.0227703
R24171 VSS.n3469 VSS.n3195 0.0227703
R24172 VSS.n4250 VSS.n2961 0.0227703
R24173 VSS.n4252 VSS.n4251 0.0227703
R24174 VSS.n2507 VSS.n2506 0.0227703
R24175 VSS.n2505 VSS.n1890 0.0227703
R24176 VSS.n2173 VSS.n2029 0.0227703
R24177 VSS.n2174 VSS.n2028 0.0227703
R24178 VSS.n218 VSS.n146 0.022693
R24179 VSS.n220 VSS.n148 0.022693
R24180 VSS.n1341 VSS.n321 0.022693
R24181 VSS.n1339 VSS.n320 0.022693
R24182 VSS.n745 VSS 0.0209651
R24183 VSS.n216 VSS.n145 0.0207632
R24184 VSS.n190 VSS.n149 0.0207632
R24185 VSS.n1343 VSS.n315 0.0207632
R24186 VSS.n1337 VSS.n317 0.0207632
R24187 VSS.n359 VSS.n358 0.0203359
R24188 VSS.n3292 VSS.n3291 0.0188784
R24189 VSS.n3300 VSS.n3299 0.0188784
R24190 VSS.n3309 VSS.n3308 0.0188784
R24191 VSS.n3318 VSS.n3317 0.0188784
R24192 VSS.n3325 VSS.n3324 0.0188784
R24193 VSS.n3351 VSS.n3350 0.0188784
R24194 VSS.n3359 VSS.n3358 0.0188784
R24195 VSS.n3368 VSS.n3367 0.0188784
R24196 VSS.n3215 VSS.n3210 0.0188784
R24197 VSS.n3443 VSS.n3211 0.0188784
R24198 VSS.n3386 VSS.n3385 0.0188784
R24199 VSS.n3418 VSS.n3391 0.0188784
R24200 VSS.n3397 VSS.n3396 0.0188784
R24201 VSS.n3400 VSS.n2931 0.0188784
R24202 VSS.n4288 VSS.n2932 0.0188784
R24203 VSS.n2941 VSS.n2940 0.0188784
R24204 VSS.n4268 VSS.n2944 0.0188784
R24205 VSS.n3951 VSS.n2946 0.0188784
R24206 VSS.n3968 VSS.n3967 0.0188784
R24207 VSS.n3928 VSS.n3927 0.0188784
R24208 VSS.n3987 VSS.n3921 0.0188784
R24209 VSS.n3990 VSS.n3989 0.0188784
R24210 VSS.n4005 VSS.n3914 0.0188784
R24211 VSS.n3705 VSS.n3080 0.0188784
R24212 VSS.n3718 VSS.n3081 0.0188784
R24213 VSS.n3710 VSS.n3075 0.0188784
R24214 VSS.n3728 VSS.n3727 0.0188784
R24215 VSS.n3733 VSS.n3732 0.0188784
R24216 VSS.n3747 VSS.n3067 0.0188784
R24217 VSS.n3745 VSS.n3061 0.0188784
R24218 VSS.n3761 VSS.n3760 0.0188784
R24219 VSS.n3766 VSS.n3765 0.0188784
R24220 VSS.n3768 VSS.n3047 0.0188784
R24221 VSS.n3775 VSS.n3048 0.0188784
R24222 VSS.n3052 VSS.n3043 0.0188784
R24223 VSS.n3786 VSS.n3783 0.0188784
R24224 VSS.n3784 VSS.n3038 0.0188784
R24225 VSS.n3799 VSS.n3039 0.0188784
R24226 VSS.n3794 VSS.n3033 0.0188784
R24227 VSS.n3811 VSS.n3810 0.0188784
R24228 VSS.n3819 VSS.n3818 0.0188784
R24229 VSS.n3827 VSS.n3021 0.0188784
R24230 VSS.n3837 VSS.n3023 0.0188784
R24231 VSS.n3845 VSS.n3017 0.0188784
R24232 VSS.n3850 VSS.n3015 0.0188784
R24233 VSS.n3853 VSS.n3852 0.0188784
R24234 VSS.n3268 VSS.n3194 0.0188784
R24235 VSS.n3472 VSS.n3471 0.0188784
R24236 VSS.n3481 VSS.n3480 0.0188784
R24237 VSS.n3483 VSS.n3185 0.0188784
R24238 VSS.n3568 VSS.n3136 0.0188784
R24239 VSS.n3580 VSS.n3138 0.0188784
R24240 VSS.n3598 VSS.n3131 0.0188784
R24241 VSS.n3590 VSS.n3132 0.0188784
R24242 VSS.n4031 VSS.n4030 0.0188784
R24243 VSS.n4040 VSS.n4039 0.0188784
R24244 VSS.n4044 VSS.n4043 0.0188784
R24245 VSS.n4048 VSS.n3895 0.0188784
R24246 VSS.n4109 VSS.n4108 0.0188784
R24247 VSS.n4113 VSS.n4112 0.0188784
R24248 VSS.n4120 VSS.n3877 0.0188784
R24249 VSS.n4123 VSS.n4122 0.0188784
R24250 VSS.n1668 VSS.n1667 0.0188784
R24251 VSS.n1672 VSS.n1671 0.0188784
R24252 VSS.n1676 VSS.n1675 0.0188784
R24253 VSS.n1680 VSS.n1679 0.0188784
R24254 VSS.n1685 VSS.n1684 0.0188784
R24255 VSS.n1697 VSS.n1696 0.0188784
R24256 VSS.n1702 VSS.n1701 0.0188784
R24257 VSS.n1705 VSS.n1704 0.0188784
R24258 VSS.n1713 VSS.n1712 0.0188784
R24259 VSS.n1717 VSS.n1716 0.0188784
R24260 VSS.n1722 VSS.n1720 0.0188784
R24261 VSS.n1731 VSS.n1730 0.0188784
R24262 VSS.n1735 VSS.n1734 0.0188784
R24263 VSS.n1739 VSS.n1738 0.0188784
R24264 VSS.n1743 VSS.n1742 0.0188784
R24265 VSS.n1748 VSS.n1747 0.0188784
R24266 VSS.n1751 VSS.n1750 0.0188784
R24267 VSS.n1759 VSS.n1758 0.0188784
R24268 VSS.n1768 VSS.n1767 0.0188784
R24269 VSS.n1778 VSS.n1777 0.0188784
R24270 VSS.n1782 VSS.n1781 0.0188784
R24271 VSS.n1786 VSS.n1785 0.0188784
R24272 VSS.n1791 VSS.n1790 0.0188784
R24273 VSS.n2205 VSS.n2204 0.0188784
R24274 VSS.n2213 VSS.n2212 0.0188784
R24275 VSS.n2222 VSS.n2221 0.0188784
R24276 VSS.n2232 VSS.n2231 0.0188784
R24277 VSS.n2241 VSS.n2240 0.0188784
R24278 VSS.n2256 VSS.n1985 0.0188784
R24279 VSS.n2277 VSS.n1987 0.0188784
R24280 VSS.n2286 VSS.n1978 0.0188784
R24281 VSS.n1980 VSS.n1975 0.0188784
R24282 VSS.n2306 VSS.n1968 0.0188784
R24283 VSS.n2309 VSS.n2308 0.0188784
R24284 VSS.n2330 VSS.n1961 0.0188784
R24285 VSS.n2339 VSS.n2338 0.0188784
R24286 VSS.n2352 VSS.n1950 0.0188784
R24287 VSS.n2354 VSS.n1941 0.0188784
R24288 VSS.n2373 VSS.n1943 0.0188784
R24289 VSS.n2386 VSS.n1936 0.0188784
R24290 VSS.n2400 VSS.n1930 0.0188784
R24291 VSS.n2417 VSS.n2416 0.0188784
R24292 VSS.n2427 VSS.n2425 0.0188784
R24293 VSS.n1913 VSS.n1907 0.0188784
R24294 VSS.n2465 VSS.n1908 0.0188784
R24295 VSS.n2443 VSS.n2442 0.0188784
R24296 VSS.n2504 VSS.n1894 0.0188784
R24297 VSS.n2494 VSS.n1889 0.0188784
R24298 VSS.n2514 VSS.n2511 0.0188784
R24299 VSS.n2512 VSS.n1883 0.0188784
R24300 VSS.n2597 VSS.n1840 0.0188784
R24301 VSS.n2603 VSS.n1841 0.0188784
R24302 VSS.n1846 VSS.n1836 0.0188784
R24303 VSS.n2613 VSS.n2611 0.0188784
R24304 VSS.n2172 VSS.n2031 0.0188784
R24305 VSS.n2163 VSS.n2055 0.0188784
R24306 VSS.n2100 VSS.n2056 0.0188784
R24307 VSS.n2104 VSS.n2103 0.0188784
R24308 VSS.n2781 VSS.n2780 0.0188784
R24309 VSS.n2777 VSS.n2776 0.0188784
R24310 VSS.n2772 VSS.n2771 0.0188784
R24311 VSS.n2768 VSS.n2767 0.0188784
R24312 VSS.n195 VSS.n144 0.0188333
R24313 VSS.n227 VSS.n150 0.0188333
R24314 VSS.n1410 VSS.n157 0.0188333
R24315 VSS.n2822 VSS.n2821 0.0188333
R24316 VSS.n1391 VSS.n296 0.0188333
R24317 VSS.n1345 VSS.n322 0.0188333
R24318 VSS.n1335 VSS.n319 0.0188333
R24319 VSS.n3276 VSS.n3275 0.0187703
R24320 VSS.n3291 VSS.n3246 0.0187703
R24321 VSS.n3336 VSS.n3334 0.0187703
R24322 VSS.n3350 VSS.n3226 0.0187703
R24323 VSS.n3389 VSS.n3386 0.0187703
R24324 VSS.n3952 VSS.n3951 0.0187703
R24325 VSS.n3960 VSS.n3959 0.0187703
R24326 VSS.n4006 VSS.n4005 0.0187703
R24327 VSS.n4015 VSS.n4014 0.0187703
R24328 VSS.n3702 VSS.n3086 0.0187703
R24329 VSS.n3705 VSS.n3704 0.0187703
R24330 VSS.n3735 VSS.n3066 0.0187703
R24331 VSS.n3751 VSS.n3067 0.0187703
R24332 VSS.n3054 VSS.n3048 0.0187703
R24333 VSS.n3820 VSS.n3819 0.0187703
R24334 VSS.n3825 VSS.n3824 0.0187703
R24335 VSS.n3853 VSS.n3009 0.0187703
R24336 VSS.n4194 VSS.n3010 0.0187703
R24337 VSS.n3497 VSS.n3181 0.0187703
R24338 VSS.n3506 VSS.n3175 0.0187703
R24339 VSS.n3508 VSS.n3172 0.0187703
R24340 VSS.n3514 VSS.n3173 0.0187703
R24341 VSS.n3533 VSS.n3532 0.0187703
R24342 VSS.n3524 VSS.n3168 0.0187703
R24343 VSS.n3527 VSS.n3525 0.0187703
R24344 VSS.n3543 VSS.n3542 0.0187703
R24345 VSS.n3545 VSS.n3153 0.0187703
R24346 VSS.n3560 VSS.n3154 0.0187703
R24347 VSS.n3551 VSS.n3149 0.0187703
R24348 VSS.n3571 VSS.n3570 0.0187703
R24349 VSS.n3607 VSS.n3122 0.0187703
R24350 VSS.n3609 VSS.n3118 0.0187703
R24351 VSS.n3621 VSS.n3119 0.0187703
R24352 VSS.n3615 VSS.n3114 0.0187703
R24353 VSS.n3634 VSS.n3633 0.0187703
R24354 VSS.n3642 VSS.n3641 0.0187703
R24355 VSS.n3647 VSS.n3646 0.0187703
R24356 VSS.n3649 VSS.n3101 0.0187703
R24357 VSS.n3670 VSS.n3102 0.0187703
R24358 VSS.n3656 VSS.n3097 0.0187703
R24359 VSS.n3680 VSS.n3678 0.0187703
R24360 VSS.n3689 VSS.n3092 0.0187703
R24361 VSS.n4054 VSS.n4053 0.0187703
R24362 VSS.n4058 VSS.n4057 0.0187703
R24363 VSS.n4063 VSS.n3891 0.0187703
R24364 VSS.n4066 VSS.n4065 0.0187703
R24365 VSS.n4069 VSS.n4068 0.0187703
R24366 VSS.n4079 VSS.n4078 0.0187703
R24367 VSS.n4083 VSS.n4082 0.0187703
R24368 VSS.n4087 VSS.n4086 0.0187703
R24369 VSS.n4091 VSS.n4090 0.0187703
R24370 VSS.n4095 VSS.n4094 0.0187703
R24371 VSS.n4102 VSS.n3881 0.0187703
R24372 VSS.n4105 VSS.n4104 0.0187703
R24373 VSS.n4130 VSS.n4129 0.0187703
R24374 VSS.n4137 VSS.n3873 0.0187703
R24375 VSS.n4140 VSS.n4139 0.0187703
R24376 VSS.n4145 VSS.n4144 0.0187703
R24377 VSS.n4148 VSS.n4147 0.0187703
R24378 VSS.n4157 VSS.n4156 0.0187703
R24379 VSS.n4161 VSS.n4160 0.0187703
R24380 VSS.n4165 VSS.n4164 0.0187703
R24381 VSS.n4169 VSS.n4168 0.0187703
R24382 VSS.n4176 VSS.n3864 0.0187703
R24383 VSS.n4179 VSS.n4178 0.0187703
R24384 VSS.n4184 VSS.n4183 0.0187703
R24385 VSS.n1663 VSS.n1662 0.0187703
R24386 VSS.n1667 VSS.n1560 0.0187703
R24387 VSS.n1688 VSS.n1687 0.0187703
R24388 VSS.n1696 VSS.n1695 0.0187703
R24389 VSS.n1722 VSS.n1721 0.0187703
R24390 VSS.n1760 VSS.n1759 0.0187703
R24391 VSS.n1765 VSS.n1764 0.0187703
R24392 VSS.n1792 VSS.n1791 0.0187703
R24393 VSS.n1797 VSS.n1795 0.0187703
R24394 VSS.n2189 VSS.n2188 0.0187703
R24395 VSS.n2204 VSS.n2018 0.0187703
R24396 VSS.n2248 VSS.n2247 0.0187703
R24397 VSS.n2256 VSS.n2255 0.0187703
R24398 VSS.n2308 VSS.n1960 0.0187703
R24399 VSS.n2401 VSS.n2400 0.0187703
R24400 VSS.n2409 VSS.n2408 0.0187703
R24401 VSS.n2443 VSS.n1903 0.0187703
R24402 VSS.n2475 VSS.n2474 0.0187703
R24403 VSS.n2522 VSS.n1879 0.0187703
R24404 VSS.n2536 VSS.n2533 0.0187703
R24405 VSS.n2534 VSS.n1869 0.0187703
R24406 VSS.n2548 VSS.n1870 0.0187703
R24407 VSS.n1873 VSS.n1865 0.0187703
R24408 VSS.n2559 VSS.n2558 0.0187703
R24409 VSS.n2564 VSS.n2563 0.0187703
R24410 VSS.n2566 VSS.n1857 0.0187703
R24411 VSS.n2579 VSS.n1858 0.0187703
R24412 VSS.n2571 VSS.n1853 0.0187703
R24413 VSS.n2590 VSS.n2589 0.0187703
R24414 VSS.n2595 VSS.n2594 0.0187703
R24415 VSS.n2626 VSS.n1831 0.0187703
R24416 VSS.n2618 VSS.n1826 0.0187703
R24417 VSS.n2637 VSS.n2636 0.0187703
R24418 VSS.n2642 VSS.n2641 0.0187703
R24419 VSS.n2644 VSS.n1819 0.0187703
R24420 VSS.n2657 VSS.n1820 0.0187703
R24421 VSS.n2653 VSS.n1815 0.0187703
R24422 VSS.n2668 VSS.n2665 0.0187703
R24423 VSS.n2666 VSS.n1810 0.0187703
R24424 VSS.n2681 VSS.n1811 0.0187703
R24425 VSS.n2676 VSS.n1806 0.0187703
R24426 VSS.n2690 VSS.n2689 0.0187703
R24427 VSS.n2116 VSS.n2115 0.0187703
R24428 VSS.n2112 VSS.n2111 0.0187703
R24429 VSS.n2125 VSS.n2124 0.0187703
R24430 VSS.n2130 VSS.n2129 0.0187703
R24431 VSS.n2134 VSS.n2133 0.0187703
R24432 VSS.n2086 VSS.n2082 0.0187703
R24433 VSS.n2084 VSS.n2069 0.0187703
R24434 VSS.n2143 VSS.n2070 0.0187703
R24435 VSS.n2075 VSS.n1449 0.0187703
R24436 VSS.n2800 VSS.n1450 0.0187703
R24437 VSS.n2793 VSS.n2792 0.0187703
R24438 VSS.n2788 VSS.n2787 0.0187703
R24439 VSS.n1586 VSS.n1469 0.0187703
R24440 VSS.n1584 VSS.n1582 0.0187703
R24441 VSS.n1595 VSS.n1594 0.0187703
R24442 VSS.n1600 VSS.n1599 0.0187703
R24443 VSS.n1608 VSS.n1607 0.0187703
R24444 VSS.n1605 VSS.n1603 0.0187703
R24445 VSS.n1618 VSS.n1617 0.0187703
R24446 VSS.n1622 VSS.n1621 0.0187703
R24447 VSS.n1629 VSS.n1628 0.0187703
R24448 VSS.n1626 VSS.n1624 0.0187703
R24449 VSS.n1642 VSS.n1641 0.0187703
R24450 VSS.n1646 VSS.n1645 0.0187703
R24451 VSS.n3299 VSS.n3199 0.0185541
R24452 VSS.n3989 VSS.n2958 0.0185541
R24453 VSS.n3719 VSS.n3718 0.0185541
R24454 VSS.n3851 VSS.n3850 0.0185541
R24455 VSS.n1671 VSS.n1492 0.0185541
R24456 VSS.n1786 VSS.n1521 0.0185541
R24457 VSS.n2212 VSS.n2014 0.0185541
R24458 VSS.n2441 VSS.n1908 0.0185541
R24459 VSS.n3489 VSS.n3186 0.0184459
R24460 VSS.n3593 VSS.n3591 0.0184459
R24461 VSS.n4050 VSS.n2968 0.0184459
R24462 VSS.n4126 VSS.n2989 0.0184459
R24463 VSS.n2525 VSS.n1884 0.0184459
R24464 VSS.n2627 VSS.n1830 0.0184459
R24465 VSS.n2106 VSS.n2060 0.0184459
R24466 VSS.n2763 VSS.n2762 0.0184459
R24467 VSS.n3391 VSS.n2928 0.0182297
R24468 VSS.n3053 VSS.n3052 0.0182297
R24469 VSS.n1730 VSS.n1506 0.0182297
R24470 VSS.n2331 VSS.n2330 0.0182297
R24471 VSS.n3490 VSS.n3489 0.0181216
R24472 VSS.n3594 VSS.n3593 0.0181216
R24473 VSS.n4050 VSS.n4049 0.0181216
R24474 VSS.n4126 VSS.n2988 0.0181216
R24475 VSS.n2526 VSS.n2525 0.0181216
R24476 VSS.n2612 VSS.n1830 0.0181216
R24477 VSS.n2106 VSS.n2059 0.0181216
R24478 VSS.n2763 VSS.n1465 0.0181216
R24479 VSS.n3336 VSS.n3335 0.0175811
R24480 VSS.n3959 VSS.n3935 0.0175811
R24481 VSS.n3752 VSS.n3066 0.0175811
R24482 VSS.n3824 VSS.n3027 0.0175811
R24483 VSS.n1687 VSS.n1553 0.0175811
R24484 VSS.n1764 VSS.n1515 0.0175811
R24485 VSS.n2248 VSS.n1994 0.0175811
R24486 VSS.n2408 VSS.n1926 0.0175811
R24487 VSS.n3497 VSS.n3496 0.0173649
R24488 VSS.n3608 VSS.n3607 0.0173649
R24489 VSS.n4054 VSS.n2969 0.0173649
R24490 VSS.n4130 VSS.n2990 0.0173649
R24491 VSS.n2532 VSS.n1879 0.0173649
R24492 VSS.n2617 VSS.n1831 0.0173649
R24493 VSS.n2116 VSS.n2061 0.0173649
R24494 VSS.n1586 VSS.n1585 0.0173649
R24495 VSS.n3483 VSS.n3482 0.0170405
R24496 VSS.n3597 VSS.n3132 0.0170405
R24497 VSS.n3895 VSS.n2965 0.0170405
R24498 VSS.n4122 VSS.n4121 0.0170405
R24499 VSS.n2513 VSS.n2512 0.0170405
R24500 VSS.n2611 VSS.n2610 0.0170405
R24501 VSS.n2103 VSS.n2097 0.0170405
R24502 VSS.n2768 VSS.n1463 0.0170405
R24503 VSS.n1420 VSS.n128 0.0169035
R24504 VSS.n229 VSS.n151 0.0169035
R24505 VSS.n276 VSS.n135 0.0169035
R24506 VSS.n1412 VSS.n156 0.0169035
R24507 VSS.n1388 VSS.n1387 0.0169035
R24508 VSS.n306 VSS.n301 0.0169035
R24509 VSS.n1347 VSS.n314 0.0169035
R24510 VSS.n1333 VSS.n318 0.0169035
R24511 VSS.n3358 VSS.n3207 0.0167162
R24512 VSS.n4268 VSS.n4267 0.0167162
R24513 VSS.n3746 VSS.n3745 0.0167162
R24514 VSS.n3810 VSS.n3029 0.0167162
R24515 VSS.n1701 VSS.n1500 0.0167162
R24516 VSS.n1750 VSS.n1540 0.0167162
R24517 VSS.n2278 VSS.n2277 0.0167162
R24518 VSS.n2386 VSS.n2385 0.0167162
R24519 VSS.n3507 VSS.n3506 0.0162838
R24520 VSS.n3622 VSS.n3118 0.0162838
R24521 VSS.n4058 VSS.n2970 0.0162838
R24522 VSS.n4138 VSS.n4137 0.0162838
R24523 VSS.n2536 VSS.n2535 0.0162838
R24524 VSS.n2635 VSS.n1826 0.0162838
R24525 VSS.n2111 VSS.n2091 0.0162838
R24526 VSS.n1582 VSS.n1475 0.0162838
R24527 VSS.n3384 VSS.n3211 0.0159595
R24528 VSS.n3400 VSS.n2927 0.0159595
R24529 VSS.n3776 VSS.n3047 0.0159595
R24530 VSS.n3785 VSS.n3784 0.0159595
R24531 VSS.n3480 VSS.n3188 0.0159595
R24532 VSS.n3137 VSS.n3131 0.0159595
R24533 VSS.n4043 VSS.n2964 0.0159595
R24534 VSS.n3877 VSS.n2985 0.0159595
R24535 VSS.n1717 VSS.n1505 0.0159595
R24536 VSS.n1738 VSS.n1544 0.0159595
R24537 VSS.n2307 VSS.n2306 0.0159595
R24538 VSS.n2337 VSS.n1950 0.0159595
R24539 VSS.n2511 VSS.n2510 0.0159595
R24540 VSS.n1846 VSS.n1845 0.0159595
R24541 VSS.n2162 VSS.n2056 0.0159595
R24542 VSS.n2772 VSS.n1445 0.0159595
R24543 VSS.n3275 VSS.n3198 0.0157432
R24544 VSS.n4014 VSS.n2959 0.0157432
R24545 VSS.n3703 VSS.n3702 0.0157432
R24546 VSS.n4195 VSS.n4194 0.0157432
R24547 VSS.n1663 VSS.n1491 0.0157432
R24548 VSS.n1795 VSS.n1522 0.0157432
R24549 VSS.n2188 VSS.n2187 0.0157432
R24550 VSS.n2475 VSS.n2472 0.0157432
R24551 VSS.n1408 VSS.n164 0.0154561
R24552 VSS.n3308 VSS.n3239 0.0152027
R24553 VSS.n3988 VSS.n3987 0.0152027
R24554 VSS.n3710 VSS.n3709 0.0152027
R24555 VSS.n3845 VSS.n3844 0.0152027
R24556 VSS.n3515 VSS.n3172 0.0152027
R24557 VSS.n3614 VSS.n3119 0.0152027
R24558 VSS.n4064 VSS.n4063 0.0152027
R24559 VSS.n4140 VSS.n2993 0.0152027
R24560 VSS.n1675 VSS.n1557 0.0152027
R24561 VSS.n1782 VSS.n1520 0.0152027
R24562 VSS.n2221 VSS.n2010 0.0152027
R24563 VSS.n2466 VSS.n1907 0.0152027
R24564 VSS.n2549 VSS.n1869 0.0152027
R24565 VSS.n2637 VSS.n1824 0.0152027
R24566 VSS.n2125 VSS.n2064 0.0152027
R24567 VSS.n1595 VSS.n1476 0.0152027
R24568 VSS.n231 VSS.n152 0.0149737
R24569 VSS.n274 VSS.n136 0.0149737
R24570 VSS.n1416 VSS.n1415 0.0149737
R24571 VSS.n1393 VSS.n295 0.0149737
R24572 VSS.n1385 VSS.n300 0.0149737
R24573 VSS.n1380 VSS.n1379 0.0149737
R24574 VSS.n1349 VSS.n323 0.0149737
R24575 VSS.n3396 VSS.n2930 0.0148784
R24576 VSS.n3783 VSS.n3782 0.0148784
R24577 VSS.n3471 VSS.n3470 0.0148784
R24578 VSS.n3581 VSS.n3580 0.0148784
R24579 VSS.n4039 VSS.n2963 0.0148784
R24580 VSS.n4112 VSS.n2984 0.0148784
R24581 VSS.n1734 VSS.n1507 0.0148784
R24582 VSS.n2339 VSS.n1956 0.0148784
R24583 VSS.n2494 VSS.n2493 0.0148784
R24584 VSS.n2604 VSS.n2603 0.0148784
R24585 VSS.n2055 VSS.n2054 0.0148784
R24586 VSS.n2777 VSS.n1447 0.0148784
R24587 VSS.n2802 VSS.n1441 0.0142297
R24588 VSS.n3324 VSS.n3204 0.0141216
R24589 VSS.n3967 VSS.n2953 0.0141216
R24590 VSS.n3734 VSS.n3733 0.0141216
R24591 VSS.n3827 VSS.n3826 0.0141216
R24592 VSS.n3173 VSS.n3166 0.0141216
R24593 VSS.n3632 VSS.n3114 0.0141216
R24594 VSS.n4066 VSS.n2973 0.0141216
R24595 VSS.n4145 VSS.n2994 0.0141216
R24596 VSS.n1685 VSS.n1497 0.0141216
R24597 VSS.n1768 VSS.n1516 0.0141216
R24598 VSS.n2241 VSS.n1998 0.0141216
R24599 VSS.n2416 VSS.n1921 0.0141216
R24600 VSS.n1872 VSS.n1870 0.0141216
R24601 VSS.n2643 VSS.n2642 0.0141216
R24602 VSS.n2130 VSS.n2065 0.0141216
R24603 VSS.n1600 VSS.n1477 0.0141216
R24604 VSS.n938 VSS.n753 0.0139402
R24605 VSS.n936 VSS.n755 0.0139402
R24606 VSS.n3693 VSS.n3692 0.0137973
R24607 VSS.n3691 VSS.n3089 0.0137973
R24608 VSS.n3569 VSS.n3568 0.0137973
R24609 VSS.n3690 VSS.n3088 0.0137973
R24610 VSS.n4108 VSS.n2983 0.0137973
R24611 VSS.n3006 VSS.n3004 0.0137973
R24612 VSS.n4201 VSS.n4200 0.0137973
R24613 VSS.n4199 VSS.n3002 0.0137973
R24614 VSS.n2698 VSS.n1524 0.0137973
R24615 VSS.n2697 VSS.n1525 0.0137973
R24616 VSS.n2597 VSS.n2596 0.0137973
R24617 VSS.n2696 VSS.n1527 0.0137973
R24618 VSS.n2780 VSS.n1444 0.0137973
R24619 VSS.n1658 VSS.n1487 0.0137973
R24620 VSS.n2743 VSS.n1488 0.0137973
R24621 VSS.n2742 VSS.n2741 0.0137973
R24622 VSS.n4187 VSS.n3859 0.0134381
R24623 VSS.n2694 VSS.n2693 0.0134381
R24624 VSS.n3367 VSS.n3208 0.0133649
R24625 VSS.n2947 VSS.n2941 0.0133649
R24626 VSS.n3760 VSS.n3759 0.0133649
R24627 VSS.n3809 VSS.n3033 0.0133649
R24628 VSS.n1705 VSS.n1501 0.0133649
R24629 VSS.n1748 VSS.n1512 0.0133649
R24630 VSS.n1986 VSS.n1978 0.0133649
R24631 VSS.n1943 VSS.n1942 0.0133649
R24632 VSS.n185 VSS.n153 0.0130439
R24633 VSS.n272 VSS.n134 0.0130439
R24634 VSS.n1377 VSS.n307 0.0130439
R24635 VSS.n1351 VSS.n313 0.0130439
R24636 VSS.n3532 VSS.n3531 0.0130405
R24637 VSS.n3633 VSS.n3110 0.0130405
R24638 VSS.n4068 VSS.n2974 0.0130405
R24639 VSS.n4147 VSS.n2995 0.0130405
R24640 VSS.n2557 VSS.n1865 0.0130405
R24641 VSS.n2658 VSS.n1819 0.0130405
R24642 VSS.n2133 VSS.n2066 0.0130405
R24643 VSS.n1607 VSS.n1606 0.0130405
R24644 VSS.n3571 VSS.n3567 0.0128243
R24645 VSS.n3679 VSS.n3092 0.0128243
R24646 VSS.n4104 VSS.n4103 0.0128243
R24647 VSS.n4183 VSS.n3003 0.0128243
R24648 VSS.n2594 VSS.n1851 0.0128243
R24649 VSS.n2690 VSS.n2688 0.0128243
R24650 VSS.n2788 VSS.n1448 0.0128243
R24651 VSS.n1646 VSS.n1486 0.0128243
R24652 VSS.n3444 VSS.n3210 0.0126081
R24653 VSS.n4289 VSS.n4288 0.0126081
R24654 VSS.n3767 VSS.n3766 0.0126081
R24655 VSS.n3800 VSS.n3799 0.0126081
R24656 VSS.n1713 VSS.n1549 0.0126081
R24657 VSS.n1742 VSS.n1510 0.0126081
R24658 VSS.n1981 VSS.n1980 0.0126081
R24659 VSS.n2354 VSS.n2353 0.0126081
R24660 VSS.n3269 VSS.n3197 0.0123919
R24661 VSS.n4028 VSS.n2960 0.0123919
R24662 VSS.n3697 VSS.n3696 0.0123919
R24663 VSS.n3861 VSS.n3860 0.0123919
R24664 VSS.n1659 VSS.n1490 0.0123919
R24665 VSS.n1796 VSS.n1526 0.0123919
R24666 VSS.n2030 VSS.n2025 0.0123919
R24667 VSS.n2473 VSS.n1893 0.0123919
R24668 VSS.n3528 VSS.n3524 0.0119595
R24669 VSS.n3642 VSS.n3107 0.0119595
R24670 VSS.n4079 VSS.n2975 0.0119595
R24671 VSS.n4157 VSS.n3869 0.0119595
R24672 VSS.n2559 VSS.n1863 0.0119595
R24673 VSS.n2652 VSS.n1820 0.0119595
R24674 VSS.n2086 VSS.n2085 0.0119595
R24675 VSS.n1603 VSS.n1480 0.0119595
R24676 VSS.n3317 VSS.n3202 0.0118514
R24677 VSS.n3927 VSS.n2955 0.0118514
R24678 VSS.n3727 VSS.n3726 0.0118514
R24679 VSS.n3023 VSS.n3022 0.0118514
R24680 VSS.n1679 VSS.n1495 0.0118514
R24681 VSS.n1778 VSS.n1536 0.0118514
R24682 VSS.n2231 VSS.n2006 0.0118514
R24683 VSS.n2427 VSS.n2426 0.0118514
R24684 VSS.n932 VSS.n931 0.01175
R24685 VSS.n929 VSS.n928 0.01175
R24686 VSS.n1146 VSS.n1145 0.01175
R24687 VSS.n1151 VSS.n1150 0.01175
R24688 VSS.n3551 VSS.n3550 0.0117432
R24689 VSS.n3678 VSS.n3677 0.0117432
R24690 VSS.n3881 VSS.n2980 0.0117432
R24691 VSS.n4178 VSS.n4177 0.0117432
R24692 VSS.n2589 VSS.n2588 0.0117432
R24693 VSS.n2676 VSS.n2675 0.0117432
R24694 VSS.n2793 VSS.n1443 0.0117432
R24695 VSS.n1641 VSS.n1485 0.0117432
R24696 VSS.n845 VSS 0.0116864
R24697 VSS.n1251 VSS 0.0116864
R24698 VSS.n3685 VSS.n3684 0.0116588
R24699 VSS.n1656 VSS.n1655 0.0116588
R24700 VSS.n3269 VSS.n3268 0.011527
R24701 VSS.n3697 VSS.n3088 0.011527
R24702 VSS.n1659 VSS.n1658 0.011527
R24703 VSS.n2172 VSS.n2030 0.011527
R24704 VSS.n4031 VSS.n4028 0.0114189
R24705 VSS.n3861 VSS.n3006 0.0114189
R24706 VSS.n2696 VSS.n1526 0.0114189
R24707 VSS.n2504 VSS.n1893 0.0114189
R24708 VSS.n238 VSS.n129 0.011114
R24709 VSS.n170 VSS.n137 0.011114
R24710 VSS VSS.n1384 0.011114
R24711 VSS.n1376 VSS.n308 0.011114
R24712 VSS.n1353 VSS.n324 0.011114
R24713 VSS.n3901 VSS.n3900 0.0109762
R24714 VSS.n3899 VSS.n3898 0.0109762
R24715 VSS.n4072 VSS.n3889 0.0109762
R24716 VSS.n4075 VSS.n4074 0.0109762
R24717 VSS.n4073 VSS.n3883 0.0109762
R24718 VSS.n4099 VSS.n4098 0.0109762
R24719 VSS.n4116 VSS.n3879 0.0109762
R24720 VSS.n4117 VSS.n3875 0.0109762
R24721 VSS.n4134 VSS.n4133 0.0109762
R24722 VSS.n4151 VSS.n3871 0.0109762
R24723 VSS.n4153 VSS.n4152 0.0109762
R24724 VSS.n4172 VSS.n3866 0.0109762
R24725 VSS.n4173 VSS.n3859 0.0109762
R24726 VSS.n3708 VSS.n3084 0.0109762
R24727 VSS.n3715 VSS.n3708 0.0109762
R24728 VSS.n3715 VSS.n3714 0.0109762
R24729 VSS.n3714 VSS.n3070 0.0109762
R24730 VSS.n3738 VSS.n3070 0.0109762
R24731 VSS.n3739 VSS.n3738 0.0109762
R24732 VSS.n3740 VSS.n3739 0.0109762
R24733 VSS.n3741 VSS.n3740 0.0109762
R24734 VSS.n3741 VSS.n3057 0.0109762
R24735 VSS.n3771 VSS.n3057 0.0109762
R24736 VSS.n3772 VSS.n3771 0.0109762
R24737 VSS.n3789 VSS.n3041 0.0109762
R24738 VSS.n3790 VSS.n3789 0.0109762
R24739 VSS.n3790 VSS.n3031 0.0109762
R24740 VSS.n3814 VSS.n3031 0.0109762
R24741 VSS.n3815 VSS.n3814 0.0109762
R24742 VSS.n3815 VSS.n3025 0.0109762
R24743 VSS.n3830 VSS.n3025 0.0109762
R24744 VSS.n3832 VSS.n3830 0.0109762
R24745 VSS.n3832 VSS.n3831 0.0109762
R24746 VSS.n3831 VSS.n3013 0.0109762
R24747 VSS.n3856 VSS.n3013 0.0109762
R24748 VSS.n4191 VSS.n3856 0.0109762
R24749 VSS.n3477 VSS.n3179 0.0109762
R24750 VSS.n3503 VSS.n3502 0.0109762
R24751 VSS.n3536 VSS.n3163 0.0109762
R24752 VSS.n3538 VSS.n3537 0.0109762
R24753 VSS.n3539 VSS.n3155 0.0109762
R24754 VSS.n3574 VSS.n3146 0.0109762
R24755 VSS.n3575 VSS.n3128 0.0109762
R24756 VSS.n3602 VSS.n3601 0.0109762
R24757 VSS.n3603 VSS.n3120 0.0109762
R24758 VSS.n3637 VSS.n3112 0.0109762
R24759 VSS.n3638 VSS.n3105 0.0109762
R24760 VSS.n2109 VSS.n2051 0.0109762
R24761 VSS.n2121 VSS.n2120 0.0109762
R24762 VSS.n2137 VSS.n2089 0.0109762
R24763 VSS.n2139 VSS.n2138 0.0109762
R24764 VSS.n2140 VSS.n1454 0.0109762
R24765 VSS.n2797 VSS.n1455 0.0109762
R24766 VSS.n2784 VSS.n1458 0.0109762
R24767 VSS.n1467 VSS.n1466 0.0109762
R24768 VSS.n1591 VSS.n1590 0.0109762
R24769 VSS.n1611 VSS.n1575 0.0109762
R24770 VSS.n1614 VSS.n1612 0.0109762
R24771 VSS.n1654 VSS.n1653 0.0109762
R24772 VSS.n1653 VSS.n1652 0.0109762
R24773 VSS.n1652 VSS.n1651 0.0109762
R24774 VSS.n1651 VSS.n1555 0.0109762
R24775 VSS.n1691 VSS.n1555 0.0109762
R24776 VSS.n1692 VSS.n1691 0.0109762
R24777 VSS.n1692 VSS.n1551 0.0109762
R24778 VSS.n1708 VSS.n1551 0.0109762
R24779 VSS.n1709 VSS.n1708 0.0109762
R24780 VSS.n1709 VSS.n1547 0.0109762
R24781 VSS.n1725 VSS.n1547 0.0109762
R24782 VSS.n1728 VSS.n1727 0.0109762
R24783 VSS.n1727 VSS.n1726 0.0109762
R24784 VSS.n1726 VSS.n1542 0.0109762
R24785 VSS.n1754 VSS.n1542 0.0109762
R24786 VSS.n1755 VSS.n1754 0.0109762
R24787 VSS.n1755 VSS.n1538 0.0109762
R24788 VSS.n1771 VSS.n1538 0.0109762
R24789 VSS.n1774 VSS.n1771 0.0109762
R24790 VSS.n1774 VSS.n1773 0.0109762
R24791 VSS.n1773 VSS.n1772 0.0109762
R24792 VSS.n1772 VSS.n1532 0.0109762
R24793 VSS.n1800 VSS.n1532 0.0109762
R24794 VSS.n2518 VSS.n2517 0.0109762
R24795 VSS.n2539 VSS.n1875 0.0109762
R24796 VSS.n2544 VSS.n2540 0.0109762
R24797 VSS.n2543 VSS.n1861 0.0109762
R24798 VSS.n2576 VSS.n2569 0.0109762
R24799 VSS.n2575 VSS.n1849 0.0109762
R24800 VSS.n2600 VSS.n2599 0.0109762
R24801 VSS.n2616 VSS.n1834 0.0109762
R24802 VSS.n2623 VSS.n2622 0.0109762
R24803 VSS.n2647 VSS.n1822 0.0109762
R24804 VSS.n2648 VSS.n1813 0.0109762
R24805 VSS.n2672 VSS.n2671 0.0109762
R24806 VSS.n2693 VSS.n1804 0.0109762
R24807 VSS.n3900 VSS.n3899 0.01095
R24808 VSS.n3898 VSS.n3889 0.01095
R24809 VSS.n4075 VSS.n4072 0.01095
R24810 VSS.n4074 VSS.n4073 0.01095
R24811 VSS.n4098 VSS.n3883 0.01095
R24812 VSS.n4099 VSS.n3879 0.01095
R24813 VSS.n4117 VSS.n4116 0.01095
R24814 VSS.n4133 VSS.n3875 0.01095
R24815 VSS.n4134 VSS.n3871 0.01095
R24816 VSS.n4153 VSS.n4151 0.01095
R24817 VSS.n4152 VSS.n3866 0.01095
R24818 VSS.n4173 VSS.n4172 0.01095
R24819 VSS.n3772 VSS.n3041 0.01095
R24820 VSS.n4191 VSS.n4190 0.01095
R24821 VSS.n3477 VSS.n3476 0.01095
R24822 VSS.n3502 VSS.n3179 0.01095
R24823 VSS.n3503 VSS.n3163 0.01095
R24824 VSS.n3537 VSS.n3536 0.01095
R24825 VSS.n3539 VSS.n3538 0.01095
R24826 VSS.n3155 VSS.n3146 0.01095
R24827 VSS.n3575 VSS.n3574 0.01095
R24828 VSS.n3601 VSS.n3128 0.01095
R24829 VSS.n3603 VSS.n3602 0.01095
R24830 VSS.n3120 VSS.n3112 0.01095
R24831 VSS.n3638 VSS.n3637 0.01095
R24832 VSS.n3652 VSS.n3105 0.01095
R24833 VSS.n2167 VSS.n2051 0.01095
R24834 VSS.n2120 VSS.n2109 0.01095
R24835 VSS.n2121 VSS.n2089 0.01095
R24836 VSS.n2138 VSS.n2137 0.01095
R24837 VSS.n2140 VSS.n2139 0.01095
R24838 VSS.n2797 VSS.n1454 0.01095
R24839 VSS.n2784 VSS.n1455 0.01095
R24840 VSS.n1466 VSS.n1458 0.01095
R24841 VSS.n1590 VSS.n1467 0.01095
R24842 VSS.n1591 VSS.n1575 0.01095
R24843 VSS.n1612 VSS.n1611 0.01095
R24844 VSS.n1614 VSS.n1613 0.01095
R24845 VSS.n1728 VSS.n1725 0.01095
R24846 VSS.n1801 VSS.n1800 0.01095
R24847 VSS.n2518 VSS.n1875 0.01095
R24848 VSS.n2540 VSS.n2539 0.01095
R24849 VSS.n2544 VSS.n2543 0.01095
R24850 VSS.n2569 VSS.n1861 0.01095
R24851 VSS.n2576 VSS.n2575 0.01095
R24852 VSS.n2599 VSS.n1849 0.01095
R24853 VSS.n2600 VSS.n1834 0.01095
R24854 VSS.n2623 VSS.n2616 0.01095
R24855 VSS.n2622 VSS.n1822 0.01095
R24856 VSS.n2648 VSS.n2647 0.01095
R24857 VSS.n2671 VSS.n1813 0.01095
R24858 VSS.n2672 VSS.n1804 0.01095
R24859 VSS.n659 VSS.n658 0.0109327
R24860 VSS.n693 VSS.n659 0.0109327
R24861 VSS.n693 VSS.n692 0.0109327
R24862 VSS.n692 VSS.n691 0.0109327
R24863 VSS.n691 VSS.n660 0.0109327
R24864 VSS.n687 VSS.n660 0.0109327
R24865 VSS.n685 VSS.n684 0.0109327
R24866 VSS.n684 VSS.n675 0.0109327
R24867 VSS.n675 VSS.n590 0.0109327
R24868 VSS.n705 VSS.n590 0.0109327
R24869 VSS.n705 VSS.n704 0.0109327
R24870 VSS.n704 VSS.n703 0.0109327
R24871 VSS.n703 VSS.n591 0.0109327
R24872 VSS.n622 VSS.n591 0.0109327
R24873 VSS.n627 VSS.n622 0.0109327
R24874 VSS.n628 VSS.n627 0.0109327
R24875 VSS.n629 VSS.n628 0.0109327
R24876 VSS.n630 VSS.n629 0.0109327
R24877 VSS.n631 VSS.n630 0.0109327
R24878 VSS.n632 VSS.n631 0.0109327
R24879 VSS.n632 VSS.n3 0.0109327
R24880 VSS.n3525 VSS.n3157 0.0108784
R24881 VSS.n3648 VSS.n3647 0.0108784
R24882 VSS.n4083 VSS.n3886 0.0108784
R24883 VSS.n4161 VSS.n2998 0.0108784
R24884 VSS.n2565 VSS.n2564 0.0108784
R24885 VSS.n2664 VSS.n1815 0.0108784
R24886 VSS.n2144 VSS.n2069 0.0108784
R24887 VSS.n1618 VSS.n1481 0.0108784
R24888 VSS.n3318 VSS.n3203 0.0107703
R24889 VSS.n3928 VSS.n2954 0.0107703
R24890 VSS.n3728 VSS.n3073 0.0107703
R24891 VSS.n3838 VSS.n3837 0.0107703
R24892 VSS.n1680 VSS.n1496 0.0107703
R24893 VSS.n1777 VSS.n1517 0.0107703
R24894 VSS.n2232 VSS.n2002 0.0107703
R24895 VSS.n2425 VSS.n1916 0.0107703
R24896 VSS.n3561 VSS.n3560 0.0106622
R24897 VSS.n3656 VSS.n3655 0.0106622
R24898 VSS.n4094 VSS.n2979 0.0106622
R24899 VSS.n3864 VSS.n3000 0.0106622
R24900 VSS.n2571 VSS.n2570 0.0106622
R24901 VSS.n2682 VSS.n2681 0.0106622
R24902 VSS.n2801 VSS.n2800 0.0106622
R24903 VSS.n1627 VSS.n1626 0.0106622
R24904 VSS.n3684 VSS.n3084 0.0106095
R24905 VSS.n1655 VSS.n1654 0.0106095
R24906 VSS.n3215 VSS.n3209 0.0100135
R24907 VSS.n2939 VSS.n2932 0.0100135
R24908 VSS.n3765 VSS.n3059 0.0100135
R24909 VSS.n3793 VSS.n3039 0.0100135
R24910 VSS.n1712 VSS.n1502 0.0100135
R24911 VSS.n1743 VSS.n1511 0.0100135
R24912 VSS.n2285 VSS.n1975 0.0100135
R24913 VSS.n2374 VSS.n1941 0.0100135
R24914 VSS.n358 VSS.n357 0.00993894
R24915 VSS.n670 VSS.n669 0.00983051
R24916 VSS.n3544 VSS.n3543 0.0097973
R24917 VSS.n3671 VSS.n3101 0.0097973
R24918 VSS.n4087 VSS.n2978 0.0097973
R24919 VSS.n4165 VSS.n2999 0.0097973
R24920 VSS.n2580 VSS.n1857 0.0097973
R24921 VSS.n2668 VSS.n2667 0.0097973
R24922 VSS.n2074 VSS.n2070 0.0097973
R24923 VSS.n1622 VSS.n1482 0.0097973
R24924 VSS.n3686 VSS.n3685 0.00967266
R24925 VSS.n1656 VSS.n1650 0.00967266
R24926 VSS.n3545 VSS.n3544 0.00958108
R24927 VSS.n3671 VSS.n3670 0.00958108
R24928 VSS.n4090 VSS.n2978 0.00958108
R24929 VSS.n4168 VSS.n2999 0.00958108
R24930 VSS.n2580 VSS.n2579 0.00958108
R24931 VSS.n2667 VSS.n2666 0.00958108
R24932 VSS.n2075 VSS.n2074 0.00958108
R24933 VSS.n1629 VSS.n1482 0.00958108
R24934 VSS.n686 VSS.n685 0.00957647
R24935 VSS.n3368 VSS.n3209 0.00925676
R24936 VSS.n2940 VSS.n2939 0.00925676
R24937 VSS.n3761 VSS.n3059 0.00925676
R24938 VSS.n3794 VSS.n3793 0.00925676
R24939 VSS.n1704 VSS.n1502 0.00925676
R24940 VSS.n1747 VSS.n1511 0.00925676
R24941 VSS.n2286 VSS.n2285 0.00925676
R24942 VSS.n2374 VSS.n2373 0.00925676
R24943 VSS.n127 VSS.n122 0.00918421
R24944 VSS.n240 VSS.n142 0.00918421
R24945 VSS.n264 VSS.n133 0.00918421
R24946 VSS.n1373 VSS.n331 0.00918421
R24947 VSS.n1355 VSS.n312 0.00918421
R24948 VSS.n1331 VSS 0.00918421
R24949 VSS.n1330 VSS.n1329 0.00918421
R24950 VSS.n4290 VSS.n2925 0.00904054
R24951 VSS.n1148 VSS.n1147 0.00885683
R24952 VSS.n1153 VSS.n1152 0.00885683
R24953 VSS.n3554 VSS.n3146 0.00880612
R24954 VSS.n2797 VSS.n1453 0.00880612
R24955 VSS.n3561 VSS.n3153 0.00871622
R24956 VSS.n3655 VSS.n3102 0.00871622
R24957 VSS.n4091 VSS.n2979 0.00871622
R24958 VSS.n4169 VSS.n3000 0.00871622
R24959 VSS.n2570 VSS.n1858 0.00871622
R24960 VSS.n2682 VSS.n1810 0.00871622
R24961 VSS.n2801 VSS.n1449 0.00871622
R24962 VSS.n1628 VSS.n1627 0.00871622
R24963 VSS.n3325 VSS.n3203 0.0085
R24964 VSS.n3968 VSS.n2954 0.0085
R24965 VSS.n3732 VSS.n3073 0.0085
R24966 VSS.n3838 VSS.n3021 0.0085
R24967 VSS.n3542 VSS.n3157 0.0085
R24968 VSS.n3649 VSS.n3648 0.0085
R24969 VSS.n4086 VSS.n3886 0.0085
R24970 VSS.n4164 VSS.n2998 0.0085
R24971 VSS.n1684 VSS.n1496 0.0085
R24972 VSS.n1767 VSS.n1517 0.0085
R24973 VSS.n2240 VSS.n2002 0.0085
R24974 VSS.n2417 VSS.n1916 0.0085
R24975 VSS.n2566 VSS.n2565 0.0085
R24976 VSS.n2665 VSS.n2664 0.0085
R24977 VSS.n2144 VSS.n2143 0.0085
R24978 VSS.n1621 VSS.n1481 0.0085
R24979 VSS.n845 VSS.n843 0.00842373
R24980 VSS.n1251 VSS.n1250 0.00842373
R24981 VSS.n1131 VSS.n1130 0.00837413
R24982 VSS.n708 VSS.n585 0.00820507
R24983 VSS.n3902 VSS.n3901 0.00809524
R24984 VSS.n2517 VSS.n1886 0.00809524
R24985 VSS.n669 VSS.n668 0.00809159
R24986 VSS.n816 VSS.n791 0.008
R24987 VSS.n812 VSS.n810 0.008
R24988 VSS.n811 VSS.n793 0.008
R24989 VSS.n806 VSS.n804 0.008
R24990 VSS.n805 VSS.n795 0.008
R24991 VSS.n800 VSS.n799 0.008
R24992 VSS.n862 VSS.n789 0.008
R24993 VSS.n890 VSS.n771 0.008
R24994 VSS.n901 VSS.n885 0.008
R24995 VSS.n892 VSS.n773 0.008
R24996 VSS.n899 VSS.n883 0.008
R24997 VSS.n894 VSS.n775 0.008
R24998 VSS.n897 VSS.n881 0.008
R24999 VSS.n896 VSS.n777 0.008
R25000 VSS.n1216 VSS.n1215 0.008
R25001 VSS.n1205 VSS.n422 0.008
R25002 VSS.n1207 VSS.n1206 0.008
R25003 VSS.n1199 VSS.n424 0.008
R25004 VSS.n1201 VSS.n1200 0.008
R25005 VSS.n1193 VSS.n426 0.008
R25006 VSS.n1195 VSS.n1194 0.008
R25007 VSS.n1192 VSS.n1191 0.008
R25008 VSS.n409 VSS.n408 0.008
R25009 VSS.n402 VSS.n368 0.008
R25010 VSS.n404 VSS.n403 0.008
R25011 VSS.n396 VSS.n370 0.008
R25012 VSS.n398 VSS.n397 0.008
R25013 VSS.n391 VSS.n372 0.008
R25014 VSS.n392 VSS.n366 0.008
R25015 VSS.n1239 VSS.n1238 0.008
R25016 VSS.n731 VSS.n717 0.00778449
R25017 VSS.n3683 VSS.n3095 0.00778095
R25018 VSS.n1649 VSS.n1564 0.00778095
R25019 VSS.n3550 VSS.n3154 0.00763514
R25020 VSS.n3677 VSS.n3097 0.00763514
R25021 VSS.n4095 VSS.n2980 0.00763514
R25022 VSS.n4177 VSS.n4176 0.00763514
R25023 VSS.n2588 VSS.n1853 0.00763514
R25024 VSS.n2675 VSS.n1811 0.00763514
R25025 VSS.n1450 VSS.n1443 0.00763514
R25026 VSS.n1624 VSS.n1485 0.00763514
R25027 VSS.n3309 VSS.n3202 0.00741892
R25028 VSS.n3921 VSS.n2955 0.00741892
R25029 VSS.n3726 VSS.n3075 0.00741892
R25030 VSS.n3022 VSS.n3017 0.00741892
R25031 VSS.n3528 VSS.n3527 0.00741892
R25032 VSS.n3646 VSS.n3107 0.00741892
R25033 VSS.n4082 VSS.n2975 0.00741892
R25034 VSS.n4160 VSS.n3869 0.00741892
R25035 VSS.n1676 VSS.n1495 0.00741892
R25036 VSS.n1781 VSS.n1536 0.00741892
R25037 VSS.n2222 VSS.n2006 0.00741892
R25038 VSS.n2426 VSS.n1913 0.00741892
R25039 VSS.n2563 VSS.n1863 0.00741892
R25040 VSS.n2653 VSS.n2652 0.00741892
R25041 VSS.n2085 VSS.n2084 0.00741892
R25042 VSS.n1617 VSS.n1480 0.00741892
R25043 VSS.n3667 VSS.n3652 0.00725714
R25044 VSS.n1613 VSS.n1569 0.00725714
R25045 VSS.n242 VSS.n130 0.00725439
R25046 VSS.n262 VSS.n138 0.00725439
R25047 VSS.n276 VSS 0.00725439
R25048 VSS.n1371 VSS.n309 0.00725439
R25049 VSS.n1357 VSS.n325 0.00725439
R25050 VSS.n839 VSS.n760 0.00716695
R25051 VSS.n1178 VSS.n1177 0.00716695
R25052 VSS.n3686 VSS.n3683 0.00707381
R25053 VSS.n1650 VSS.n1649 0.00707381
R25054 VSS.n3276 VSS.n3197 0.00698649
R25055 VSS.n4015 VSS.n2960 0.00698649
R25056 VSS.n3696 VSS.n3086 0.00698649
R25057 VSS.n3860 VSS.n3010 0.00698649
R25058 VSS.n1662 VSS.n1490 0.00698649
R25059 VSS.n1797 VSS.n1796 0.00698649
R25060 VSS.n2189 VSS.n2025 0.00698649
R25061 VSS.n2474 VSS.n2473 0.00698649
R25062 VSS.n3476 VSS.n3192 0.00696162
R25063 VSS.n2168 VSS.n2167 0.00696162
R25064 VSS.n4190 VSS.n3857 0.00691667
R25065 VSS.n1801 VSS.n1531 0.00691667
R25066 VSS VSS.n730 0.00686346
R25067 VSS.n3444 VSS.n3443 0.00666216
R25068 VSS.n4289 VSS.n2931 0.00666216
R25069 VSS.n3768 VSS.n3767 0.00666216
R25070 VSS.n3800 VSS.n3038 0.00666216
R25071 VSS.n1716 VSS.n1549 0.00666216
R25072 VSS.n1739 VSS.n1510 0.00666216
R25073 VSS.n1981 VSS.n1968 0.00666216
R25074 VSS.n2353 VSS.n2352 0.00666216
R25075 VSS.n3567 VSS.n3149 0.00655405
R25076 VSS.n3680 VSS.n3679 0.00655405
R25077 VSS.n4103 VSS.n4102 0.00655405
R25078 VSS.n4179 VSS.n3003 0.00655405
R25079 VSS.n2590 VSS.n1851 0.00655405
R25080 VSS.n2688 VSS.n1806 0.00655405
R25081 VSS.n2792 VSS.n1448 0.00655405
R25082 VSS.n1642 VSS.n1486 0.00655405
R25083 VSS.n3531 VSS.n3168 0.00633784
R25084 VSS.n3641 VSS.n3110 0.00633784
R25085 VSS.n4078 VSS.n2974 0.00633784
R25086 VSS.n4156 VSS.n2995 0.00633784
R25087 VSS.n2558 VSS.n2557 0.00633784
R25088 VSS.n2658 VSS.n2657 0.00633784
R25089 VSS.n2082 VSS.n2066 0.00633784
R25090 VSS.n1606 VSS.n1605 0.00633784
R25091 VSS.n674 VSS.n673 0.00625916
R25092 VSS.n3359 VSS.n3208 0.00590541
R25093 VSS.n2947 VSS.n2944 0.00590541
R25094 VSS.n3759 VSS.n3061 0.00590541
R25095 VSS.n3811 VSS.n3809 0.00590541
R25096 VSS.n1702 VSS.n1501 0.00590541
R25097 VSS.n1751 VSS.n1512 0.00590541
R25098 VSS.n1987 VSS.n1986 0.00590541
R25099 VSS.n1942 VSS.n1936 0.00590541
R25100 VSS.n3141 VSS.n3128 0.00588776
R25101 VSS.n3476 VSS.n3191 0.00588776
R25102 VSS.n1461 VSS.n1458 0.00588776
R25103 VSS.n2167 VSS.n2050 0.00588776
R25104 VSS VSS.n4295 0.00555747
R25105 VSS.n3570 VSS.n3569 0.00547297
R25106 VSS.n3690 VSS.n3689 0.00547297
R25107 VSS.n4105 VSS.n2983 0.00547297
R25108 VSS.n4184 VSS.n3004 0.00547297
R25109 VSS.n2596 VSS.n2595 0.00547297
R25110 VSS.n2689 VSS.n1527 0.00547297
R25111 VSS.n2787 VSS.n1444 0.00547297
R25112 VSS.n1645 VSS.n1487 0.00547297
R25113 VSS.n180 VSS.n141 0.00532456
R25114 VSS.n260 VSS.n132 0.00532456
R25115 VSS.n1410 VSS 0.00532456
R25116 VSS.n1369 VSS.n330 0.00532456
R25117 VSS.n1359 VSS.n311 0.00532456
R25118 VSS.n3533 VSS.n3166 0.00525676
R25119 VSS.n3634 VSS.n3632 0.00525676
R25120 VSS.n4069 VSS.n2973 0.00525676
R25121 VSS.n4148 VSS.n2994 0.00525676
R25122 VSS.n1873 VSS.n1872 0.00525676
R25123 VSS.n2644 VSS.n2643 0.00525676
R25124 VSS.n2134 VSS.n2065 0.00525676
R25125 VSS.n1608 VSS.n1477 0.00525676
R25126 VSS.n3334 VSS.n3204 0.00514865
R25127 VSS.n3960 VSS.n2953 0.00514865
R25128 VSS.n4290 VSS.n2926 0.00514865
R25129 VSS.n3735 VSS.n3734 0.00514865
R25130 VSS.n3826 VSS.n3825 0.00514865
R25131 VSS.n1688 VSS.n1497 0.00514865
R25132 VSS.n1765 VSS.n1516 0.00514865
R25133 VSS.n2247 VSS.n1998 0.00514865
R25134 VSS.n2409 VSS.n1921 0.00514865
R25135 VSS.n4188 VSS.n4187 0.00440238
R25136 VSS.n2694 VSS.n1803 0.00440238
R25137 VSS.n3418 VSS.n2930 0.00439189
R25138 VSS.n3782 VSS.n3043 0.00439189
R25139 VSS.n3470 VSS.n3194 0.00439189
R25140 VSS.n3581 VSS.n3136 0.00439189
R25141 VSS.n4030 VSS.n2963 0.00439189
R25142 VSS.n4109 VSS.n2984 0.00439189
R25143 VSS.n1731 VSS.n1507 0.00439189
R25144 VSS.n1961 VSS.n1956 0.00439189
R25145 VSS.n2493 VSS.n1894 0.00439189
R25146 VSS.n2604 VSS.n1840 0.00439189
R25147 VSS.n2054 VSS.n2031 0.00439189
R25148 VSS.n2781 VSS.n1447 0.00439189
R25149 VSS.n3699 VSS.n3698 0.00425921
R25150 VSS.n3701 VSS.n3085 0.00425921
R25151 VSS.n3729 VSS.n3074 0.00425921
R25152 VSS.n3731 VSS.n3071 0.00425921
R25153 VSS.n3749 VSS.n3748 0.00425921
R25154 VSS.n3744 VSS.n3743 0.00425921
R25155 VSS.n3762 VSS.n3060 0.00425921
R25156 VSS.n3764 VSS.n3058 0.00425921
R25157 VSS.n3051 VSS.n3050 0.00425921
R25158 VSS.n3798 VSS.n3797 0.00425921
R25159 VSS.n3795 VSS.n3032 0.00425921
R25160 VSS.n3812 VSS.n3030 0.00425921
R25161 VSS.n3817 VSS.n3028 0.00425921
R25162 VSS.n3828 VSS.n3024 0.00425921
R25163 VSS.n3836 VSS.n3835 0.00425921
R25164 VSS.n4193 VSS.n3011 0.00425921
R25165 VSS.n3862 VSS.n3012 0.00425921
R25166 VSS.n3541 VSS.n3158 0.00425921
R25167 VSS.n3546 VSS.n3156 0.00425921
R25168 VSS.n3650 VSS.n3106 0.00425921
R25169 VSS.n3669 VSS.n3103 0.00425921
R25170 VSS.n4047 VSS.n4046 0.00425921
R25171 VSS.n4052 VSS.n4051 0.00425921
R25172 VSS.n4056 VSS.n4055 0.00425921
R25173 VSS.n4060 VSS.n4059 0.00425921
R25174 VSS.n4081 VSS.n4080 0.00425921
R25175 VSS.n4085 VSS.n4084 0.00425921
R25176 VSS.n4089 VSS.n4088 0.00425921
R25177 VSS.n4093 VSS.n4092 0.00425921
R25178 VSS.n4110 VSS.n4107 0.00425921
R25179 VSS.n4124 VSS.n3876 0.00425921
R25180 VSS.n4128 VSS.n4127 0.00425921
R25181 VSS.n4131 VSS.n3874 0.00425921
R25182 VSS.n4136 VSS.n3872 0.00425921
R25183 VSS.n4159 VSS.n4158 0.00425921
R25184 VSS.n4163 VSS.n4162 0.00425921
R25185 VSS.n4167 VSS.n4166 0.00425921
R25186 VSS.n4170 VSS.n3865 0.00425921
R25187 VSS.n1661 VSS.n1660 0.00425921
R25188 VSS.n1665 VSS.n1664 0.00425921
R25189 VSS.n1681 VSS.n1678 0.00425921
R25190 VSS.n1686 VSS.n1683 0.00425921
R25191 VSS.n1698 VSS.n1552 0.00425921
R25192 VSS.n1703 VSS.n1700 0.00425921
R25193 VSS.n1706 VSS.n1550 0.00425921
R25194 VSS.n1714 VSS.n1711 0.00425921
R25195 VSS.n1732 VSS.n1729 0.00425921
R25196 VSS.n1744 VSS.n1741 0.00425921
R25197 VSS.n1749 VSS.n1746 0.00425921
R25198 VSS.n1752 VSS.n1541 0.00425921
R25199 VSS.n1757 VSS.n1539 0.00425921
R25200 VSS.n1769 VSS.n1537 0.00425921
R25201 VSS.n1779 VSS.n1776 0.00425921
R25202 VSS.n1794 VSS.n1793 0.00425921
R25203 VSS.n1798 VSS.n1528 0.00425921
R25204 VSS.n1888 VSS.n1885 0.00425921
R25205 VSS.n2524 VSS.n2523 0.00425921
R25206 VSS.n2520 VSS.n1876 0.00425921
R25207 VSS.n2537 VSS.n1878 0.00425921
R25208 VSS.n2562 VSS.n2560 0.00425921
R25209 VSS.n2567 VSS.n1862 0.00425921
R25210 VSS.n2578 VSS.n1859 0.00425921
R25211 VSS.n2572 VSS.n1860 0.00425921
R25212 VSS.n2598 VSS.n1842 0.00425921
R25213 VSS.n2614 VSS.n1835 0.00425921
R25214 VSS.n2625 VSS.n1832 0.00425921
R25215 VSS.n2619 VSS.n1833 0.00425921
R25216 VSS.n2620 VSS.n1825 0.00425921
R25217 VSS.n2655 VSS.n2654 0.00425921
R25218 VSS.n2650 VSS.n1814 0.00425921
R25219 VSS.n2669 VSS.n1812 0.00425921
R25220 VSS.n2680 VSS.n2674 0.00425921
R25221 VSS.n2142 VSS.n2071 0.00425921
R25222 VSS.n2077 VSS.n2076 0.00425921
R25223 VSS.n1620 VSS.n1619 0.00425921
R25224 VSS.n1630 VSS.n1623 0.00425921
R25225 VSS.n3665 VSS.n3664 0.00424524
R25226 VSS.n1635 VSS.n1634 0.00424524
R25227 VSS.n3706 VSS.n3085 0.0042371
R25228 VSS.n3717 VSS.n3082 0.0042371
R25229 VSS.n3711 VSS.n3083 0.0042371
R25230 VSS.n3712 VSS.n3074 0.0042371
R25231 VSS.n3736 VSS.n3072 0.0042371
R25232 VSS.n3750 VSS.n3749 0.0042371
R25233 VSS.n3769 VSS.n3058 0.0042371
R25234 VSS.n3774 VSS.n3049 0.0042371
R25235 VSS.n3056 VSS.n3055 0.0042371
R25236 VSS.n3055 VSS.n3051 0.0042371
R25237 VSS.n3050 VSS.n3042 0.0042371
R25238 VSS.n3787 VSS.n3040 0.0042371
R25239 VSS.n3798 VSS.n3792 0.0042371
R25240 VSS.n3821 VSS.n3028 0.0042371
R25241 VSS.n3823 VSS.n3026 0.0042371
R25242 VSS.n3835 VSS.n3834 0.0042371
R25243 VSS.n3847 VSS.n3846 0.0042371
R25244 VSS.n3849 VSS.n3014 0.0042371
R25245 VSS.n3854 VSS.n3011 0.0042371
R25246 VSS.n3484 VSS.n3187 0.0042371
R25247 VSS.n3513 VSS.n3164 0.0042371
R25248 VSS.n3534 VSS.n3165 0.0042371
R25249 VSS.n3572 VSS.n3148 0.0042371
R25250 VSS.n3599 VSS.n3130 0.0042371
R25251 VSS.n3616 VSS.n3113 0.0042371
R25252 VSS.n3635 VSS.n3111 0.0042371
R25253 VSS.n3681 VSS.n3096 0.0042371
R25254 VSS.n3688 VSS.n3093 0.0042371
R25255 VSS.n4042 VSS.n4041 0.0042371
R25256 VSS.n4046 VSS.n4045 0.0042371
R25257 VSS.n4062 VSS.n4060 0.0042371
R25258 VSS.n4067 VSS.n3890 0.0042371
R25259 VSS.n4070 VSS.n3888 0.0042371
R25260 VSS.n4080 VSS.n4077 0.0042371
R25261 VSS.n4096 VSS.n4093 0.0042371
R25262 VSS.n4101 VSS.n3882 0.0042371
R25263 VSS.n4106 VSS.n3880 0.0042371
R25264 VSS.n4107 VSS.n4106 0.0042371
R25265 VSS.n4111 VSS.n4110 0.0042371
R25266 VSS.n4114 VSS.n3878 0.0042371
R25267 VSS.n4119 VSS.n3876 0.0042371
R25268 VSS.n4141 VSS.n3872 0.0042371
R25269 VSS.n4146 VSS.n4143 0.0042371
R25270 VSS.n4149 VSS.n3870 0.0042371
R25271 VSS.n4158 VSS.n4155 0.0042371
R25272 VSS.n4175 VSS.n3865 0.0042371
R25273 VSS.n4180 VSS.n3863 0.0042371
R25274 VSS.n4185 VSS.n4182 0.0042371
R25275 VSS.n4186 VSS.n4185 0.0042371
R25276 VSS.n1666 VSS.n1665 0.0042371
R25277 VSS.n1670 VSS.n1669 0.0042371
R25278 VSS.n1674 VSS.n1673 0.0042371
R25279 VSS.n1678 VSS.n1677 0.0042371
R25280 VSS.n1689 VSS.n1554 0.0042371
R25281 VSS.n1694 VSS.n1552 0.0042371
R25282 VSS.n1715 VSS.n1714 0.0042371
R25283 VSS.n1719 VSS.n1718 0.0042371
R25284 VSS.n1723 VSS.n1546 0.0042371
R25285 VSS.n1729 VSS.n1546 0.0042371
R25286 VSS.n1733 VSS.n1732 0.0042371
R25287 VSS.n1737 VSS.n1736 0.0042371
R25288 VSS.n1741 VSS.n1740 0.0042371
R25289 VSS.n1761 VSS.n1539 0.0042371
R25290 VSS.n1766 VSS.n1763 0.0042371
R25291 VSS.n1780 VSS.n1779 0.0042371
R25292 VSS.n1784 VSS.n1783 0.0042371
R25293 VSS.n1789 VSS.n1787 0.0042371
R25294 VSS.n1793 VSS.n1533 0.0042371
R25295 VSS.n2496 VSS.n1887 0.0042371
R25296 VSS.n2515 VSS.n1888 0.0042371
R25297 VSS.n1878 VSS.n1877 0.0042371
R25298 VSS.n2547 VSS.n2546 0.0042371
R25299 VSS.n2541 VSS.n1874 0.0042371
R25300 VSS.n2560 VSS.n1864 0.0042371
R25301 VSS.n2573 VSS.n2572 0.0042371
R25302 VSS.n2591 VSS.n1852 0.0042371
R25303 VSS.n2593 VSS.n1850 0.0042371
R25304 VSS.n2598 VSS.n1850 0.0042371
R25305 VSS.n2602 VSS.n1842 0.0042371
R25306 VSS.n1848 VSS.n1847 0.0042371
R25307 VSS.n1843 VSS.n1835 0.0042371
R25308 VSS.n2638 VSS.n1825 0.0042371
R25309 VSS.n2640 VSS.n1823 0.0042371
R25310 VSS.n2645 VSS.n1821 0.0042371
R25311 VSS.n2656 VSS.n2655 0.0042371
R25312 VSS.n2680 VSS.n2679 0.0042371
R25313 VSS.n2677 VSS.n1805 0.0042371
R25314 VSS.n2691 VSS.n1529 0.0042371
R25315 VSS.n2695 VSS.n1529 0.0042371
R25316 VSS.n2102 VSS.n2101 0.0042371
R25317 VSS.n2131 VSS.n2128 0.0042371
R25318 VSS.n2135 VSS.n2132 0.0042371
R25319 VSS.n2789 VSS.n2786 0.0042371
R25320 VSS.n2770 VSS.n2769 0.0042371
R25321 VSS.n1601 VSS.n1598 0.0042371
R25322 VSS.n1609 VSS.n1602 0.0042371
R25323 VSS.n1643 VSS.n1640 0.0042371
R25324 VSS.n1647 VSS.n1644 0.0042371
R25325 VSS.n4034 VSS.n4033 0.00423273
R25326 VSS.n2502 VSS.n2501 0.00423273
R25327 VSS.n2786 VSS.n2785 0.00423268
R25328 VSS.n3264 VSS.n3263 0.00422178
R25329 VSS.n4021 VSS.n3905 0.00422178
R25330 VSS.n2490 VSS.n2489 0.00422178
R25331 VSS.n2045 VSS.n2044 0.00422178
R25332 VSS.n3667 VSS.n3666 0.00421905
R25333 VSS.n1633 VSS.n1569 0.00421905
R25334 VSS.n3515 VSS.n3514 0.00417568
R25335 VSS.n3615 VSS.n3614 0.00417568
R25336 VSS.n4065 VSS.n4064 0.00417568
R25337 VSS.n4144 VSS.n2993 0.00417568
R25338 VSS.n2549 VSS.n2548 0.00417568
R25339 VSS.n2641 VSS.n1824 0.00417568
R25340 VSS.n2129 VSS.n2064 0.00417568
R25341 VSS.n1599 VSS.n1476 0.00417568
R25342 VSS.n3707 VSS.n3082 0.00410442
R25343 VSS.n3855 VSS.n3014 0.00410442
R25344 VSS.n1669 VSS.n1559 0.00410442
R25345 VSS.n1789 VSS.n1788 0.00410442
R25346 VSS.n3300 VSS.n3239 0.00406757
R25347 VSS.n3990 VSS.n3988 0.00406757
R25348 VSS.n3709 VSS.n3081 0.00406757
R25349 VSS.n3844 VSS.n3015 0.00406757
R25350 VSS.n1672 VSS.n1557 0.00406757
R25351 VSS.n1785 VSS.n1520 0.00406757
R25352 VSS.n2213 VSS.n2010 0.00406757
R25353 VSS.n2466 VSS.n2465 0.00406757
R25354 VSS.n3553 VSS.n3147 0.00402269
R25355 VSS.n2791 VSS.n1456 0.00402269
R25356 VSS.n3488 VSS.n3177 0.00398793
R25357 VSS.n3592 VSS.n3125 0.00398793
R25358 VSS.n2107 VSS.n2094 0.00398793
R25359 VSS.n2764 VSS.n1468 0.00398793
R25360 VSS.n4051 VSS.n3894 0.00397174
R25361 VSS.n4089 VSS.n3884 0.00397174
R25362 VSS.n4127 VSS.n4125 0.00397174
R25363 VSS.n4171 VSS.n4167 0.00397174
R25364 VSS.n2524 VSS.n2519 0.00397174
R25365 VSS.n2578 VSS.n2577 0.00397174
R25366 VSS.n2615 VSS.n1832 0.00397174
R25367 VSS.n2673 VSS.n1812 0.00397174
R25368 VSS.n2802 VSS.n1442 0.00395946
R25369 VSS.n3763 VSS.n3762 0.00394963
R25370 VSS.n3796 VSS.n3795 0.00394963
R25371 VSS.n1710 VSS.n1550 0.00394963
R25372 VSS.n1746 VSS.n1745 0.00394963
R25373 VSS.n3479 VSS.n3189 0.00394626
R25374 VSS.n3140 VSS.n3129 0.00394626
R25375 VSS.n2098 VSS.n2053 0.00394626
R25376 VSS.n2774 VSS.n2773 0.00394626
R25377 VSS.n3256 VSS.n3190 0.00393696
R25378 VSS.n3578 VSS.n3577 0.00393696
R25379 VSS.n2049 VSS.n2048 0.00393696
R25380 VSS.n2782 VSS.n2779 0.00393696
R25381 VSS.n3498 VSS.n3176 0.00390294
R25382 VSS.n3610 VSS.n3121 0.00390294
R25383 VSS.n2114 VSS.n2113 0.00390294
R25384 VSS.n1583 VSS.n1581 0.00390294
R25385 VSS.n3559 VSS.n3558 0.00389381
R25386 VSS.n2799 VSS.n2798 0.00389381
R25387 VSS.n3509 VSS.n3174 0.00385851
R25388 VSS.n3523 VSS.n3159 0.00385851
R25389 VSS.n3620 VSS.n3613 0.00385851
R25390 VSS.n3644 VSS.n3643 0.00385851
R25391 VSS.n2123 VSS.n2122 0.00385851
R25392 VSS.n2087 VSS.n2078 0.00385851
R25393 VSS.n1593 VSS.n1592 0.00385851
R25394 VSS.n1615 VSS.n1572 0.00385851
R25395 VSS.n3510 VSS.n3509 0.00380768
R25396 VSS.n3620 VSS.n3619 0.00380768
R25397 VSS.n2123 VSS.n2090 0.00380768
R25398 VSS.n1593 VSS.n1576 0.00380768
R25399 VSS.n3523 VSS.n3162 0.00380053
R25400 VSS.n3643 VSS.n3109 0.00380053
R25401 VSS.n2088 VSS.n2087 0.00380053
R25402 VSS.n1574 VSS.n1572 0.00380053
R25403 VSS.n3731 VSS.n3730 0.00379484
R25404 VSS.n3833 VSS.n3024 0.00379484
R25405 VSS.n4032 VSS.n3904 0.00379484
R25406 VSS.n1683 VSS.n1682 0.00379484
R25407 VSS.n1775 VSS.n1537 0.00379484
R25408 VSS.n2503 VSS.n1897 0.00379484
R25409 VSS.n3687 VSS.n3094 0.00377273
R25410 VSS.n1657 VSS.n1563 0.00377273
R25411 VSS.n3485 VSS.n3484 0.0037725
R25412 VSS.n3559 VSS.n3549 0.0037725
R25413 VSS.n3130 VSS.n3126 0.0037725
R25414 VSS.n2102 VSS.n2096 0.0037725
R25415 VSS.n2799 VSS.n1451 0.0037725
R25416 VSS.n2769 VSS.n1464 0.0037725
R25417 VSS.n3663 VSS.n3662 0.00374762
R25418 VSS.n1637 VSS.n1636 0.00374762
R25419 VSS.n3577 VSS.n3576 0.00372958
R25420 VSS.n4061 VSS.n3890 0.0037285
R25421 VSS.n4143 VSS.n4142 0.0037285
R25422 VSS.n2547 VSS.n1871 0.0037285
R25423 VSS.n2640 VSS.n2639 0.0037285
R25424 VSS.n3148 VSS.n3145 0.00372177
R25425 VSS.n4076 VSS.n3888 0.00370639
R25426 VSS.n4154 VSS.n3870 0.00370639
R25427 VSS.n2542 VSS.n2541 0.00370639
R25428 VSS.n2649 VSS.n1821 0.00370639
R25429 VSS.n3661 VSS.n3095 0.00369524
R25430 VSS.n1638 VSS.n1564 0.00369524
R25431 VSS.n3072 VSS.n3068 0.00366216
R25432 VSS.n3823 VSS.n3822 0.00366216
R25433 VSS.n3654 VSS.n3653 0.00366216
R25434 VSS.n1693 VSS.n1554 0.00366216
R25435 VSS.n1763 VSS.n1762 0.00366216
R25436 VSS.n1568 VSS.n1567 0.00366216
R25437 VSS.n3668 VSS.n3104 0.00364005
R25438 VSS.n1632 VSS.n1631 0.00364005
R25439 VSS.n3246 VSS.n3198 0.00363514
R25440 VSS.n4006 VSS.n2959 0.00363514
R25441 VSS.n3704 VSS.n3703 0.00363514
R25442 VSS.n4195 VSS.n3009 0.00363514
R25443 VSS.n1560 VSS.n1491 0.00363514
R25444 VSS.n1792 VSS.n1522 0.00363514
R25445 VSS.n2187 VSS.n2018 0.00363514
R25446 VSS.n2472 VSS.n1903 0.00363514
R25447 VSS.n1131 VSS.n1113 0.00362312
R25448 VSS.n4037 VSS.n4035 0.00359048
R25449 VSS.n2500 VSS.n2499 0.00359048
R25450 VSS.n3547 VSS.n3546 0.00358532
R25451 VSS.n2076 VSS.n2073 0.00358532
R25452 VSS.n2783 VSS.n1457 0.00358218
R25453 VSS.n3263 VSS.n3259 0.00357902
R25454 VSS.n4021 VSS.n4020 0.00357902
R25455 VSS.n2044 VSS.n2034 0.00357902
R25456 VSS.n2489 VSS.n1898 0.00357902
R25457 VSS.n3488 VSS.n3487 0.00357098
R25458 VSS.n3592 VSS.n3127 0.00357098
R25459 VSS.n2108 VSS.n2107 0.00357098
R25460 VSS.n2765 VSS.n2764 0.00357098
R25461 VSS.n3744 VSS.n3069 0.00348526
R25462 VSS.n3816 VSS.n3030 0.00348526
R25463 VSS.n1700 VSS.n1699 0.00348526
R25464 VSS.n1756 VSS.n1541 0.00348526
R25465 VSS.n3513 VSS.n3512 0.003457
R25466 VSS.n3617 VSS.n3616 0.003457
R25467 VSS.n2128 VSS.n2127 0.003457
R25468 VSS.n1598 VSS.n1597 0.003457
R25469 VSS.n3165 VSS.n3161 0.00344926
R25470 VSS.n3639 VSS.n3111 0.00344926
R25471 VSS.n2132 VSS.n2080 0.00344926
R25472 VSS.n1602 VSS.n1573 0.00344926
R25473 VSS.n4056 VSS.n3892 0.00344103
R25474 VSS.n4084 VSS.n3887 0.00344103
R25475 VSS.n4135 VSS.n3874 0.00344103
R25476 VSS.n4162 VSS.n3868 0.00344103
R25477 VSS.n2538 VSS.n1876 0.00344103
R25478 VSS.n2561 VSS.n1862 0.00344103
R25479 VSS.n2621 VSS.n2619 0.00344103
R25480 VSS.n2651 VSS.n2650 0.00344103
R25481 VSS.n3526 VSS.n3160 0.00343273
R25482 VSS.n3645 VSS.n3108 0.00343273
R25483 VSS.n2083 VSS.n2079 0.00343273
R25484 VSS.n1616 VSS.n1571 0.00343273
R25485 VSS.n3505 VSS.n3504 0.00341839
R25486 VSS.n3612 VSS.n3611 0.00341839
R25487 VSS.n2093 VSS.n2092 0.00341839
R25488 VSS.n1578 VSS.n1577 0.00341839
R25489 VSS.n3604 VSS.n3603 0.00341837
R25490 VSS.n3502 VSS.n3178 0.00341837
R25491 VSS.n1590 VSS.n1579 0.00341837
R25492 VSS.n2120 VSS.n2095 0.00341837
R25493 VSS.n249 VSS.n131 0.00339474
R25494 VSS.n175 VSS.n139 0.00339474
R25495 VSS.n1367 VSS.n310 0.00339474
R25496 VSS.n1361 VSS.n328 0.00339474
R25497 VSS.n4036 VSS.n3902 0.00335476
R25498 VSS.n2498 VSS.n1886 0.00335476
R25499 VSS.n3713 VSS.n3711 0.00335258
R25500 VSS.n3846 VSS.n3016 0.00335258
R25501 VSS.n1674 VSS.n1556 0.00335258
R25502 VSS.n1783 VSS.n1535 0.00335258
R25503 VSS.n3504 VSS.n3176 0.0033136
R25504 VSS.n3611 VSS.n3610 0.0033136
R25505 VSS.n2113 VSS.n2093 0.0033136
R25506 VSS.n1583 VSS.n1578 0.0033136
R25507 VSS.n3385 VSS.n3384 0.00331081
R25508 VSS.n3397 VSS.n2927 0.00331081
R25509 VSS.n3776 VSS.n3775 0.00331081
R25510 VSS.n3786 VSS.n3785 0.00331081
R25511 VSS.n3472 VSS.n3188 0.00331081
R25512 VSS.n3138 VSS.n3137 0.00331081
R25513 VSS.n4040 VSS.n2964 0.00331081
R25514 VSS.n4113 VSS.n2985 0.00331081
R25515 VSS.n1720 VSS.n1505 0.00331081
R25516 VSS.n1735 VSS.n1544 0.00331081
R25517 VSS.n2309 VSS.n2307 0.00331081
R25518 VSS.n2338 VSS.n2337 0.00331081
R25519 VSS.n2510 VSS.n1889 0.00331081
R25520 VSS.n1845 VSS.n1841 0.00331081
R25521 VSS.n2163 VSS.n2162 0.00331081
R25522 VSS.n2776 VSS.n1445 0.00331081
R25523 VSS.n3167 VSS.n3161 0.00330444
R25524 VSS.n3640 VSS.n3639 0.00330444
R25525 VSS.n2081 VSS.n2080 0.00330444
R25526 VSS.n1604 VSS.n1573 0.00330444
R25527 VSS.n3160 VSS.n3158 0.0032992
R25528 VSS.n3108 VSS.n3106 0.0032992
R25529 VSS.n2079 VSS.n2071 0.0032992
R25530 VSS.n1619 VSS.n1571 0.0032992
R25531 VSS.n3512 VSS.n3511 0.00329663
R25532 VSS.n3618 VSS.n3617 0.00329663
R25533 VSS.n2127 VSS.n2126 0.00329663
R25534 VSS.n1597 VSS.n1596 0.00329663
R25535 VSS.n3659 VSS.n3658 0.00324201
R25536 VSS.n1566 VSS.n1565 0.00324201
R25537 VSS.n3770 VSS.n3049 0.00319779
R25538 VSS.n3791 VSS.n3040 0.00319779
R25539 VSS.n3660 VSS.n3096 0.00319779
R25540 VSS.n4097 VSS.n3882 0.00319779
R25541 VSS.n4174 VSS.n3863 0.00319779
R25542 VSS.n1718 VSS.n1548 0.00319779
R25543 VSS.n1737 VSS.n1543 0.00319779
R25544 VSS.n2574 VSS.n1852 0.00319779
R25545 VSS.n2678 VSS.n2677 0.00319779
R25546 VSS.n1640 VSS.n1639 0.00319779
R25547 VSS.n3479 VSS.n3478 0.00317568
R25548 VSS.n3600 VSS.n3129 0.00317568
R25549 VSS.n4042 VSS.n3896 0.00317568
R25550 VSS.n4118 VSS.n3878 0.00317568
R25551 VSS.n2516 VSS.n1887 0.00317568
R25552 VSS.n1847 VSS.n1844 0.00317568
R25553 VSS.n2099 VSS.n2098 0.00317568
R25554 VSS.n2773 VSS.n1462 0.00317568
R25555 VSS.n3487 VSS.n3486 0.00316007
R25556 VSS.n3589 VSS.n3127 0.00316007
R25557 VSS.n2108 VSS.n2105 0.00316007
R25558 VSS.n2766 VSS.n2765 0.00316007
R25559 VSS.n3548 VSS.n3547 0.00314581
R25560 VSS.n2073 VSS.n2072 0.00314581
R25561 VSS.n4038 VSS.n3903 0.00310934
R25562 VSS.n2495 VSS.n2492 0.00310934
R25563 VSS.n3508 VSS.n3507 0.00309459
R25564 VSS.n3622 VSS.n3621 0.00309459
R25565 VSS.n3891 VSS.n2970 0.00309459
R25566 VSS.n4139 VSS.n4138 0.00309459
R25567 VSS.n2535 VSS.n2534 0.00309459
R25568 VSS.n2636 VSS.n2635 0.00309459
R25569 VSS.n2124 VSS.n2091 0.00309459
R25570 VSS.n1594 VSS.n1475 0.00309459
R25571 VSS.n3700 VSS.n3699 0.003043
R25572 VSS.n4192 VSS.n3012 0.003043
R25573 VSS.n1661 VSS.n1561 0.003043
R25574 VSS.n1799 VSS.n1798 0.003043
R25575 VSS.n3576 VSS.n3144 0.00302306
R25576 VSS.n3145 VSS.n3144 0.00300884
R25577 VSS.n3305 VSS.n3303 0.0029881
R25578 VSS.n3340 VSS.n3339 0.0029881
R25579 VSS.n3355 VSS.n3221 0.0029881
R25580 VSS.n3941 VSS.n2943 0.0029881
R25581 VSS.n2218 VSS.n2216 0.0029881
R25582 VSS.n2251 VSS.n1996 0.0029881
R25583 VSS.n2274 VSS.n2266 0.0029881
R25584 VSS.n2390 VSS.n2389 0.0029881
R25585 VSS.n3549 VSS.n3548 0.00298054
R25586 VSS.n3486 VSS.n3485 0.00298054
R25587 VSS.n3589 VSS.n3126 0.00298054
R25588 VSS.n2105 VSS.n2096 0.00298054
R25589 VSS.n2072 VSS.n1451 0.00298054
R25590 VSS.n2766 VSS.n1464 0.00298054
R25591 VSS.n3956 VSS.n3933 0.0029619
R25592 VSS.n3985 VSS.n3984 0.0029619
R25593 VSS.n2405 VSS.n1924 0.0029619
R25594 VSS.n2437 VSS.n2436 0.0029619
R25595 VSS.n3167 VSS.n3162 0.00293083
R25596 VSS.n3640 VSS.n3109 0.00293083
R25597 VSS.n2088 VSS.n2081 0.00293083
R25598 VSS.n1604 VSS.n1574 0.00293083
R25599 VSS.n3511 VSS.n3510 0.0029237
R25600 VSS.n3619 VSS.n3618 0.0029237
R25601 VSS.n2126 VSS.n2090 0.0029237
R25602 VSS.n1596 VSS.n1576 0.0029237
R25603 VSS.n3774 VSS.n3773 0.00291032
R25604 VSS.n3788 VSS.n3787 0.00291032
R25605 VSS.n3573 VSS.n3147 0.00291032
R25606 VSS.n3682 VSS.n3681 0.00291032
R25607 VSS.n4041 VSS.n3897 0.00291032
R25608 VSS.n4101 VSS.n4100 0.00291032
R25609 VSS.n4115 VSS.n4114 0.00291032
R25610 VSS.n4181 VSS.n4180 0.00291032
R25611 VSS.n1724 VSS.n1719 0.00291032
R25612 VSS.n1736 VSS.n1545 0.00291032
R25613 VSS.n2497 VSS.n2496 0.00291032
R25614 VSS.n2592 VSS.n2591 0.00291032
R25615 VSS.n2601 VSS.n1848 0.00291032
R25616 VSS.n2692 VSS.n1805 0.00291032
R25617 VSS.n2791 VSS.n2790 0.00291032
R25618 VSS.n1648 VSS.n1643 0.00291032
R25619 VSS.n3505 VSS.n3174 0.00289527
R25620 VSS.n3613 VSS.n3612 0.00289527
R25621 VSS.n3526 VSS.n3159 0.00289527
R25622 VSS.n3645 VSS.n3644 0.00289527
R25623 VSS.n2122 VSS.n2092 0.00289527
R25624 VSS.n2083 VSS.n2078 0.00289527
R25625 VSS.n1592 VSS.n1577 0.00289527
R25626 VSS.n1616 VSS.n1615 0.00289527
R25627 VSS.n3261 VSS.n3259 0.00287188
R25628 VSS.n2042 VSS.n2034 0.00287188
R25629 VSS.n4023 VSS.n4020 0.00284569
R25630 VSS.n2487 VSS.n1898 0.00284569
R25631 VSS.n3558 VSS.n3557 0.00283826
R25632 VSS.n2798 VSS.n1452 0.00283826
R25633 VSS.n4188 VSS.n3857 0.00283095
R25634 VSS.n1803 VSS.n1531 0.00283095
R25635 VSS.n3193 VSS.n3190 0.00279542
R25636 VSS.n3579 VSS.n3578 0.00279542
R25637 VSS.n2052 VSS.n2049 0.00279542
R25638 VSS.n2779 VSS.n2778 0.00279542
R25639 VSS.n3180 VSS.n3177 0.00276679
R25640 VSS.n3125 VSS.n3124 0.00276679
R25641 VSS.n2110 VSS.n2094 0.00276679
R25642 VSS.n1580 VSS.n1468 0.00276679
R25643 VSS.n3716 VSS.n3083 0.00275553
R25644 VSS.n3848 VSS.n3847 0.00275553
R25645 VSS.n1673 VSS.n1558 0.00275553
R25646 VSS.n1784 VSS.n1534 0.00275553
R25647 VSS.n488 VSS.n487 0.00274058
R25648 VSS.n1023 VSS.n479 0.00274058
R25649 VSS.n1043 VSS.n471 0.00274058
R25650 VSS.n1064 VSS.n1060 0.00274058
R25651 VSS.n3698 VSS.n3087 0.00273342
R25652 VSS.n4186 VSS.n3862 0.00273342
R25653 VSS.n1660 VSS.n1562 0.00273342
R25654 VSS.n2695 VSS.n1528 0.00273342
R25655 VSS.n3261 VSS.n3260 0.00272619
R25656 VSS.n3260 VSS.n3253 0.00272619
R25657 VSS.n3279 VSS.n3251 0.00272619
R25658 VSS.n3281 VSS.n3280 0.00272619
R25659 VSS.n3289 VSS.n3288 0.00272619
R25660 VSS.n3297 VSS.n3241 0.00272619
R25661 VSS.n3302 VSS.n3241 0.00272619
R25662 VSS.n3304 VSS.n3237 0.00272619
R25663 VSS.n3312 VSS.n3237 0.00272619
R25664 VSS.n3320 VSS.n3234 0.00272619
R25665 VSS.n3321 VSS.n3320 0.00272619
R25666 VSS.n3330 VSS.n3329 0.00272619
R25667 VSS.n3331 VSS.n3330 0.00272619
R25668 VSS.n3341 VSS.n3228 0.00272619
R25669 VSS.n3345 VSS.n3228 0.00272619
R25670 VSS.n3353 VSS.n3224 0.00272619
R25671 VSS.n3354 VSS.n3353 0.00272619
R25672 VSS.n3362 VSS.n3361 0.00272619
R25673 VSS.n3365 VSS.n3364 0.00272619
R25674 VSS.n3374 VSS.n3373 0.00272619
R25675 VSS.n3441 VSS.n3440 0.00272619
R25676 VSS.n3440 VSS.n3439 0.00272619
R25677 VSS.n3434 VSS.n3433 0.00272619
R25678 VSS.n3433 VSS.n3383 0.00272619
R25679 VSS.n3429 VSS.n3383 0.00272619
R25680 VSS.n3423 VSS.n3422 0.00272619
R25681 VSS.n3414 VSS.n3413 0.00272619
R25682 VSS.n3413 VSS.n3395 0.00272619
R25683 VSS.n3407 VSS.n3399 0.00272619
R25684 VSS.n3403 VSS.n3399 0.00272619
R25685 VSS.n3403 VSS.n3402 0.00272619
R25686 VSS.n4284 VSS.n4283 0.00272619
R25687 VSS.n4283 VSS.n2936 0.00272619
R25688 VSS.n4274 VSS.n2938 0.00272619
R25689 VSS.n4274 VSS.n4273 0.00272619
R25690 VSS.n3946 VSS.n3940 0.00272619
R25691 VSS.n3955 VSS.n3954 0.00272619
R25692 VSS.n3963 VSS.n3962 0.00272619
R25693 VSS.n3965 VSS.n3964 0.00272619
R25694 VSS.n3973 VSS.n3925 0.00272619
R25695 VSS.n3983 VSS.n3982 0.00272619
R25696 VSS.n3985 VSS.n3983 0.00272619
R25697 VSS.n3993 VSS.n3919 0.00272619
R25698 VSS.n3994 VSS.n3993 0.00272619
R25699 VSS.n3995 VSS.n3994 0.00272619
R25700 VSS.n4003 VSS.n4001 0.00272619
R25701 VSS.n4003 VSS.n4002 0.00272619
R25702 VSS.n4012 VSS.n4010 0.00272619
R25703 VSS.n4012 VSS.n4011 0.00272619
R25704 VSS.n4026 VSS.n4025 0.00272619
R25705 VSS.n4024 VSS.n4023 0.00272619
R25706 VSS.n2042 VSS.n2041 0.00272619
R25707 VSS.n2041 VSS.n2040 0.00272619
R25708 VSS.n2192 VSS.n2023 0.00272619
R25709 VSS.n2194 VSS.n2193 0.00272619
R25710 VSS.n2202 VSS.n2201 0.00272619
R25711 VSS.n2210 VSS.n2012 0.00272619
R25712 VSS.n2215 VSS.n2012 0.00272619
R25713 VSS.n2217 VSS.n2008 0.00272619
R25714 VSS.n2225 VSS.n2008 0.00272619
R25715 VSS.n2227 VSS.n2004 0.00272619
R25716 VSS.n2235 VSS.n2004 0.00272619
R25717 VSS.n2243 VSS.n2000 0.00272619
R25718 VSS.n2244 VSS.n2243 0.00272619
R25719 VSS.n2253 VSS.n2252 0.00272619
R25720 VSS.n2253 VSS.n1992 0.00272619
R25721 VSS.n2261 VSS.n1990 0.00272619
R25722 VSS.n2265 VSS.n1990 0.00272619
R25723 VSS.n2273 VSS.n2272 0.00272619
R25724 VSS.n2268 VSS.n2267 0.00272619
R25725 VSS.n2291 VSS.n1973 0.00272619
R25726 VSS.n2301 VSS.n2300 0.00272619
R25727 VSS.n2304 VSS.n2301 0.00272619
R25728 VSS.n2312 VSS.n1966 0.00272619
R25729 VSS.n2313 VSS.n2312 0.00272619
R25730 VSS.n2314 VSS.n2313 0.00272619
R25731 VSS.n2328 VSS.n2327 0.00272619
R25732 VSS.n2342 VSS.n1954 0.00272619
R25733 VSS.n2343 VSS.n2342 0.00272619
R25734 VSS.n2349 VSS.n2348 0.00272619
R25735 VSS.n2350 VSS.n2349 0.00272619
R25736 VSS.n2350 VSS.n1948 0.00272619
R25737 VSS.n2359 VSS.n1946 0.00272619
R25738 VSS.n2363 VSS.n1946 0.00272619
R25739 VSS.n2369 VSS.n2368 0.00272619
R25740 VSS.n2368 VSS.n2365 0.00272619
R25741 VSS.n2395 VSS.n1932 0.00272619
R25742 VSS.n2404 VSS.n2403 0.00272619
R25743 VSS.n2412 VSS.n2411 0.00272619
R25744 VSS.n2414 VSS.n2413 0.00272619
R25745 VSS.n2423 VSS.n2422 0.00272619
R25746 VSS.n2432 VSS.n1911 0.00272619
R25747 VSS.n2436 VSS.n1911 0.00272619
R25748 VSS.n2463 VSS.n2462 0.00272619
R25749 VSS.n2462 VSS.n2461 0.00272619
R25750 VSS.n2461 VSS.n2438 0.00272619
R25751 VSS.n2452 VSS.n2440 0.00272619
R25752 VSS.n2452 VSS.n2451 0.00272619
R25753 VSS.n2445 VSS.n1901 0.00272619
R25754 VSS.n2478 VSS.n1901 0.00272619
R25755 VSS.n2485 VSS.n2484 0.00272619
R25756 VSS.n2487 VSS.n2486 0.00272619
R25757 VSS.n3271 VSS.n3253 0.0027
R25758 VSS.n3280 VSS.n3279 0.0027
R25759 VSS.n3289 VSS.n3287 0.0027
R25760 VSS.n3297 VSS.n3296 0.0027
R25761 VSS.n3305 VSS.n3304 0.0027
R25762 VSS.n3331 VSS.n3230 0.0027
R25763 VSS.n3365 VSS.n3362 0.0027
R25764 VSS.n3373 VSS.n3372 0.0027
R25765 VSS.n3441 VSS.n3380 0.0027
R25766 VSS.n3423 VSS.n3388 0.0027
R25767 VSS.n3415 VSS.n3414 0.0027
R25768 VSS.n4273 VSS.n4272 0.0027
R25769 VSS.n3942 VSS.n3940 0.0027
R25770 VSS.n3954 VSS.n3937 0.0027
R25771 VSS.n3965 VSS.n3963 0.0027
R25772 VSS.n3973 VSS.n3972 0.0027
R25773 VSS.n3982 VSS.n3923 0.0027
R25774 VSS.n4011 VSS.n3909 0.0027
R25775 VSS.n4025 VSS.n4024 0.0027
R25776 VSS.n2040 VSS.n2039 0.0027
R25777 VSS.n2193 VSS.n2192 0.0027
R25778 VSS.n2202 VSS.n2200 0.0027
R25779 VSS.n2210 VSS.n2209 0.0027
R25780 VSS.n2218 VSS.n2217 0.0027
R25781 VSS.n2245 VSS.n2244 0.0027
R25782 VSS.n2272 VSS.n2267 0.0027
R25783 VSS.n2291 VSS.n2290 0.0027
R25784 VSS.n2300 VSS.n1971 0.0027
R25785 VSS.n2328 VSS.n2320 0.0027
R25786 VSS.n2321 VSS.n1954 0.0027
R25787 VSS.n2365 VSS.n1934 0.0027
R25788 VSS.n2391 VSS.n1932 0.0027
R25789 VSS.n2403 VSS.n1928 0.0027
R25790 VSS.n2414 VSS.n2412 0.0027
R25791 VSS.n2423 VSS.n2421 0.0027
R25792 VSS.n2432 VSS.n2431 0.0027
R25793 VSS.n2479 VSS.n2478 0.0027
R25794 VSS.n2486 VSS.n2485 0.0027
R25795 VSS.n3339 VSS.n3230 0.00264762
R25796 VSS.n3962 VSS.n3933 0.00264762
R25797 VSS.n2245 VSS.n1996 0.00264762
R25798 VSS.n2411 VSS.n1924 0.00264762
R25799 VSS.n4055 VSS.n3893 0.00264496
R25800 VSS.n4132 VSS.n4131 0.00264496
R25801 VSS.n2521 VSS.n2520 0.00264496
R25802 VSS.n2624 VSS.n1833 0.00264496
R25803 VSS.n3541 VSS.n3540 0.00262285
R25804 VSS.n3651 VSS.n3650 0.00262285
R25805 VSS.n4085 VSS.n3885 0.00262285
R25806 VSS.n4163 VSS.n3867 0.00262285
R25807 VSS.n2568 VSS.n2567 0.00262285
R25808 VSS.n2670 VSS.n1814 0.00262285
R25809 VSS.n2142 VSS.n2141 0.00262285
R25810 VSS.n1620 VSS.n1570 0.00262285
R25811 VSS.n3355 VSS.n3354 0.00262143
R25812 VSS.n3942 VSS.n3941 0.00262143
R25813 VSS.n2266 VSS.n2265 0.00262143
R25814 VSS.n2391 VSS.n2390 0.00262143
R25815 VSS.n3743 VSS.n3742 0.00260074
R25816 VSS.n3813 VSS.n3812 0.00260074
R25817 VSS.n1707 VSS.n1703 0.00260074
R25818 VSS.n1753 VSS.n1752 0.00260074
R25819 VSS.n3307 VSS.n3240 0.00257862
R25820 VSS.n3986 VSS.n3920 0.00257862
R25821 VSS.n2220 VSS.n2011 0.00257862
R25822 VSS.n2435 VSS.n1909 0.00257862
R25823 VSS.n4272 VSS.n2943 0.00256905
R25824 VSS.n2389 VSS.n1934 0.00256905
R25825 VSS.n3351 VSS.n3207 0.00255405
R25826 VSS.n4267 VSS.n2946 0.00255405
R25827 VSS.n3747 VSS.n3746 0.00255405
R25828 VSS.n3818 VSS.n3029 0.00255405
R25829 VSS.n1697 VSS.n1500 0.00255405
R25830 VSS.n1758 VSS.n1540 0.00255405
R25831 VSS.n2278 VSS.n1985 0.00255405
R25832 VSS.n2385 VSS.n1930 0.00255405
R25833 VSS.n3361 VSS.n3221 0.00254286
R25834 VSS.n3956 VSS.n3955 0.00254286
R25835 VSS.n2274 VSS.n2273 0.00254286
R25836 VSS.n2405 VSS.n2404 0.00254286
R25837 VSS.n3357 VSS.n3222 0.0025344
R25838 VSS.n2276 VSS.n2275 0.0025344
R25839 VSS.n720 VSS.n716 0.00252206
R25840 VSS.n723 VSS.n722 0.00252206
R25841 VSS.n726 VSS.n719 0.00252206
R25842 VSS.n728 VSS.n727 0.00252206
R25843 VSS.n732 VSS.n715 0.00252206
R25844 VSS.n3341 VSS.n3340 0.00251667
R25845 VSS.n2252 VSS.n2251 0.00251667
R25846 VSS.n4270 VSS.n4269 0.00251228
R25847 VSS.n2388 VSS.n2387 0.00251228
R25848 VSS.n2785 VSS.n1457 0.00249519
R25849 VSS.n3266 VSS.n3265 0.0024936
R25850 VSS.n2169 VSS.n2046 0.0024936
R25851 VSS.n3303 VSS.n3302 0.00246429
R25852 VSS.n3984 VSS.n3919 0.00246429
R25853 VSS.n2216 VSS.n2215 0.00246429
R25854 VSS.n2463 VSS.n2437 0.00246429
R25855 VSS.n3737 VSS.n3736 0.00244595
R25856 VSS.n3829 VSS.n3026 0.00244595
R25857 VSS.n1690 VSS.n1689 0.00244595
R25858 VSS.n1770 VSS.n1766 0.00244595
R25859 VSS.n3322 VSS.n3321 0.0024381
R25860 VSS.n3972 VSS.n3971 0.0024381
R25861 VSS.n2236 VSS.n2235 0.0024381
R25862 VSS.n2421 VSS.n2420 0.0024381
R25863 VSS.n3338 VSS.n3337 0.00242383
R25864 VSS.n3958 VSS.n3934 0.00242383
R25865 VSS.n2249 VSS.n1997 0.00242383
R25866 VSS.n2407 VSS.n1925 0.00242383
R25867 VSS.n4035 VSS.n4034 0.00238571
R25868 VSS.n3664 VSS.n3663 0.00238571
R25869 VSS.n3286 VSS.n3249 0.00238571
R25870 VSS.n3295 VSS.n3244 0.00238571
R25871 VSS.n3314 VSS.n3313 0.00238571
R25872 VSS.n3322 VSS.n3232 0.00238571
R25873 VSS.n3347 VSS.n3346 0.00238571
R25874 VSS.n3363 VSS.n3217 0.00238571
R25875 VSS.n3379 VSS.n3214 0.00238571
R25876 VSS.n3428 VSS.n3427 0.00238571
R25877 VSS.n3421 VSS.n3393 0.00238571
R25878 VSS.n3409 VSS.n3395 0.00238571
R25879 VSS.n4285 VSS.n2935 0.00238571
R25880 VSS.n4279 VSS.n4278 0.00238571
R25881 VSS.n3948 VSS.n3947 0.00238571
R25882 VSS.n3971 VSS.n3929 0.00238571
R25883 VSS.n3978 VSS.n3977 0.00238571
R25884 VSS.n4000 VSS.n3917 0.00238571
R25885 VSS.n4009 VSS.n3912 0.00238571
R25886 VSS.n1636 VSS.n1635 0.00238571
R25887 VSS.n2501 VSS.n2500 0.00238571
R25888 VSS.n2199 VSS.n2021 0.00238571
R25889 VSS.n2208 VSS.n2016 0.00238571
R25890 VSS.n2228 VSS.n2226 0.00238571
R25891 VSS.n2237 VSS.n2236 0.00238571
R25892 VSS.n2260 VSS.n2259 0.00238571
R25893 VSS.n2289 VSS.n1976 0.00238571
R25894 VSS.n2296 VSS.n2295 0.00238571
R25895 VSS.n2319 VSS.n1964 0.00238571
R25896 VSS.n2326 VSS.n2322 0.00238571
R25897 VSS.n2344 VSS.n2343 0.00238571
R25898 VSS.n2358 VSS.n2357 0.00238571
R25899 VSS.n2370 VSS.n2364 0.00238571
R25900 VSS.n2397 VSS.n2396 0.00238571
R25901 VSS.n2420 VSS.n1919 0.00238571
R25902 VSS.n2430 VSS.n1914 0.00238571
R25903 VSS.n2457 VSS.n2456 0.00238571
R25904 VSS.n2450 VSS.n2446 0.00238571
R25905 VSS.n3278 VSS.n3277 0.00237961
R25906 VSS.n3282 VSS.n3250 0.00237961
R25907 VSS.n3290 VSS.n3248 0.00237961
R25908 VSS.n3298 VSS.n3242 0.00237961
R25909 VSS.n3301 VSS.n3242 0.00237961
R25910 VSS.n3310 VSS.n3238 0.00237961
R25911 VSS.n3311 VSS.n3310 0.00237961
R25912 VSS.n3319 VSS.n3235 0.00237961
R25913 VSS.n3319 VSS.n3233 0.00237961
R25914 VSS.n3328 VSS.n3231 0.00237961
R25915 VSS.n3332 VSS.n3231 0.00237961
R25916 VSS.n3343 VSS.n3342 0.00237961
R25917 VSS.n3344 VSS.n3343 0.00237961
R25918 VSS.n3352 VSS.n3225 0.00237961
R25919 VSS.n3352 VSS.n3223 0.00237961
R25920 VSS.n3360 VSS.n3219 0.00237961
R25921 VSS.n3366 VSS.n3220 0.00237961
R25922 VSS.n3375 VSS.n3216 0.00237961
R25923 VSS.n3442 VSS.n3213 0.00237961
R25924 VSS.n3438 VSS.n3213 0.00237961
R25925 VSS.n3432 VSS.n3382 0.00237961
R25926 VSS.n3432 VSS.n3431 0.00237961
R25927 VSS.n3431 VSS.n3430 0.00237961
R25928 VSS.n3424 VSS.n3392 0.00237961
R25929 VSS.n3412 VSS.n3394 0.00237961
R25930 VSS.n3412 VSS.n3411 0.00237961
R25931 VSS.n3406 VSS.n3405 0.00237961
R25932 VSS.n3405 VSS.n3404 0.00237961
R25933 VSS.n3404 VSS.n3401 0.00237961
R25934 VSS.n4282 VSS.n2934 0.00237961
R25935 VSS.n4282 VSS.n4281 0.00237961
R25936 VSS.n4276 VSS.n4275 0.00237961
R25937 VSS.n4275 VSS.n2942 0.00237961
R25938 VSS.n3945 VSS.n3944 0.00237961
R25939 VSS.n3953 VSS.n3936 0.00237961
R25940 VSS.n3961 VSS.n3931 0.00237961
R25941 VSS.n3966 VSS.n3932 0.00237961
R25942 VSS.n3975 VSS.n3974 0.00237961
R25943 VSS.n3981 VSS.n3922 0.00237961
R25944 VSS.n3986 VSS.n3922 0.00237961
R25945 VSS.n3992 VSS.n3991 0.00237961
R25946 VSS.n3992 VSS.n3918 0.00237961
R25947 VSS.n3996 VSS.n3918 0.00237961
R25948 VSS.n4004 VSS.n3915 0.00237961
R25949 VSS.n4004 VSS.n3916 0.00237961
R25950 VSS.n4013 VSS.n3911 0.00237961
R25951 VSS.n4013 VSS.n3910 0.00237961
R25952 VSS.n4027 VSS.n3906 0.00237961
R25953 VSS.n3267 VSS.n3258 0.00237961
R25954 VSS.n3474 VSS.n3473 0.00237961
R25955 VSS.n3535 VSS.n3164 0.00237961
R25956 VSS.n3535 VSS.n3534 0.00237961
R25957 VSS.n3555 VSS.n3552 0.00237961
R25958 VSS.n3142 VSS.n3139 0.00237961
R25959 VSS.n3636 VSS.n3113 0.00237961
R25960 VSS.n3636 VSS.n3635 0.00237961
R25961 VSS.n4071 VSS.n4067 0.00237961
R25962 VSS.n4071 VSS.n4070 0.00237961
R25963 VSS.n4150 VSS.n4146 0.00237961
R25964 VSS.n4150 VSS.n4149 0.00237961
R25965 VSS.n2191 VSS.n2190 0.00237961
R25966 VSS.n2195 VSS.n2022 0.00237961
R25967 VSS.n2203 VSS.n2020 0.00237961
R25968 VSS.n2211 VSS.n2013 0.00237961
R25969 VSS.n2214 VSS.n2013 0.00237961
R25970 VSS.n2223 VSS.n2009 0.00237961
R25971 VSS.n2224 VSS.n2223 0.00237961
R25972 VSS.n2233 VSS.n2005 0.00237961
R25973 VSS.n2234 VSS.n2233 0.00237961
R25974 VSS.n2242 VSS.n2001 0.00237961
R25975 VSS.n2242 VSS.n1999 0.00237961
R25976 VSS.n2254 VSS.n1995 0.00237961
R25977 VSS.n2254 VSS.n1993 0.00237961
R25978 VSS.n2263 VSS.n2262 0.00237961
R25979 VSS.n2264 VSS.n2263 0.00237961
R25980 VSS.n2271 VSS.n1989 0.00237961
R25981 VSS.n2270 VSS.n2269 0.00237961
R25982 VSS.n2293 VSS.n2292 0.00237961
R25983 VSS.n2299 VSS.n1969 0.00237961
R25984 VSS.n2305 VSS.n1969 0.00237961
R25985 VSS.n2311 VSS.n2310 0.00237961
R25986 VSS.n2311 VSS.n1965 0.00237961
R25987 VSS.n2315 VSS.n1965 0.00237961
R25988 VSS.n2329 VSS.n1963 0.00237961
R25989 VSS.n2341 VSS.n2340 0.00237961
R25990 VSS.n2341 VSS.n1953 0.00237961
R25991 VSS.n2347 VSS.n1951 0.00237961
R25992 VSS.n2351 VSS.n1951 0.00237961
R25993 VSS.n2351 VSS.n1949 0.00237961
R25994 VSS.n2361 VSS.n2360 0.00237961
R25995 VSS.n2362 VSS.n2361 0.00237961
R25996 VSS.n2367 VSS.n1945 0.00237961
R25997 VSS.n2367 VSS.n2366 0.00237961
R25998 VSS.n2394 VSS.n2393 0.00237961
R25999 VSS.n2402 VSS.n1927 0.00237961
R26000 VSS.n2410 VSS.n1922 0.00237961
R26001 VSS.n2415 VSS.n1923 0.00237961
R26002 VSS.n2424 VSS.n1918 0.00237961
R26003 VSS.n2434 VSS.n2433 0.00237961
R26004 VSS.n2435 VSS.n2434 0.00237961
R26005 VSS.n2464 VSS.n1910 0.00237961
R26006 VSS.n2460 VSS.n1910 0.00237961
R26007 VSS.n2460 VSS.n2459 0.00237961
R26008 VSS.n2454 VSS.n2453 0.00237961
R26009 VSS.n2453 VSS.n2444 0.00237961
R26010 VSS.n2476 VSS.n1902 0.00237961
R26011 VSS.n2477 VSS.n2476 0.00237961
R26012 VSS.n2483 VSS.n1895 0.00237961
R26013 VSS.n2546 VSS.n2545 0.00237961
R26014 VSS.n2545 VSS.n1874 0.00237961
R26015 VSS.n2646 VSS.n1823 0.00237961
R26016 VSS.n2646 VSS.n2645 0.00237961
R26017 VSS.n2171 VSS.n2170 0.00237961
R26018 VSS.n2165 VSS.n2164 0.00237961
R26019 VSS.n2136 VSS.n2131 0.00237961
R26020 VSS.n2136 VSS.n2135 0.00237961
R26021 VSS.n2795 VSS.n2794 0.00237961
R26022 VSS.n2775 VSS.n1460 0.00237961
R26023 VSS.n1610 VSS.n1601 0.00237961
R26024 VSS.n1610 VSS.n1609 0.00237961
R26025 VSS.n3372 VSS.n3217 0.00235952
R26026 VSS.n3435 VSS.n3434 0.00235952
R26027 VSS.n2290 VSS.n2289 0.00235952
R26028 VSS.n2302 VSS.n1966 0.00235952
R26029 VSS.n3270 VSS.n3254 0.00235749
R26030 VSS.n3278 VSS.n3250 0.00235749
R26031 VSS.n3290 VSS.n3247 0.00235749
R26032 VSS.n3298 VSS.n3243 0.00235749
R26033 VSS.n3306 VSS.n3238 0.00235749
R26034 VSS.n3333 VSS.n3332 0.00235749
R26035 VSS.n3366 VSS.n3219 0.00235749
R26036 VSS.n3371 VSS.n3216 0.00235749
R26037 VSS.n3442 VSS.n3212 0.00235749
R26038 VSS.n3425 VSS.n3424 0.00235749
R26039 VSS.n3416 VSS.n3394 0.00235749
R26040 VSS.n4271 VSS.n2942 0.00235749
R26041 VSS.n3944 VSS.n3943 0.00235749
R26042 VSS.n3953 VSS.n3938 0.00235749
R26043 VSS.n3966 VSS.n3931 0.00235749
R26044 VSS.n3974 VSS.n3926 0.00235749
R26045 VSS.n3981 VSS.n3980 0.00235749
R26046 VSS.n4016 VSS.n3910 0.00235749
R26047 VSS.n3500 VSS.n3499 0.00235749
R26048 VSS.n3606 VSS.n3605 0.00235749
R26049 VSS.n2038 VSS.n2032 0.00235749
R26050 VSS.n2191 VSS.n2022 0.00235749
R26051 VSS.n2203 VSS.n2019 0.00235749
R26052 VSS.n2211 VSS.n2015 0.00235749
R26053 VSS.n2219 VSS.n2009 0.00235749
R26054 VSS.n2246 VSS.n1999 0.00235749
R26055 VSS.n2271 VSS.n2270 0.00235749
R26056 VSS.n2292 VSS.n1974 0.00235749
R26057 VSS.n2299 VSS.n2298 0.00235749
R26058 VSS.n2329 VSS.n1962 0.00235749
R26059 VSS.n2340 VSS.n1955 0.00235749
R26060 VSS.n2366 VSS.n1935 0.00235749
R26061 VSS.n2393 VSS.n2392 0.00235749
R26062 VSS.n2402 VSS.n1929 0.00235749
R26063 VSS.n2415 VSS.n1922 0.00235749
R26064 VSS.n2424 VSS.n1917 0.00235749
R26065 VSS.n2433 VSS.n1912 0.00235749
R26066 VSS.n2477 VSS.n1900 0.00235749
R26067 VSS.n2118 VSS.n2117 0.00235749
R26068 VSS.n1588 VSS.n1587 0.00235749
R26069 VSS.n4279 VSS.n2936 0.00233333
R26070 VSS.n2364 VSS.n2363 0.00233333
R26071 VSS.n3338 VSS.n3333 0.00231327
R26072 VSS.n3961 VSS.n3934 0.00231327
R26073 VSS.n2246 VSS.n1997 0.00231327
R26074 VSS.n2410 VSS.n1925 0.00231327
R26075 VSS.n3272 VSS.n3271 0.00230714
R26076 VSS.n4018 VSS.n3909 0.00230714
R26077 VSS.n4026 VSS.n4019 0.00230714
R26078 VSS.n2039 VSS.n2036 0.00230714
R26079 VSS.n2480 VSS.n2479 0.00230714
R26080 VSS.n2484 VSS.n1899 0.00230714
R26081 VSS.n3356 VSS.n3223 0.00229115
R26082 VSS.n3943 VSS.n2945 0.00229115
R26083 VSS.n3737 VSS.n3071 0.00229115
R26084 VSS.n3829 VSS.n3828 0.00229115
R26085 VSS.n1690 VSS.n1686 0.00229115
R26086 VSS.n1770 VSS.n1769 0.00229115
R26087 VSS.n2264 VSS.n1988 0.00229115
R26088 VSS.n2392 VSS.n1933 0.00229115
R26089 VSS.n3273 VSS.n3251 0.00228095
R26090 VSS.n3288 VSS.n3244 0.00228095
R26091 VSS.n2035 VSS.n2023 0.00228095
R26092 VSS.n2201 VSS.n2016 0.00228095
R26093 VSS.n4001 VSS.n4000 0.00225476
R26094 VSS.n2456 VSS.n2440 0.00225476
R26095 VSS.n4271 VSS.n4270 0.00224693
R26096 VSS.n2388 VSS.n1935 0.00224693
R26097 VSS.n3482 VSS.n3481 0.00222973
R26098 VSS.n3598 VSS.n3597 0.00222973
R26099 VSS.n4044 VSS.n2965 0.00222973
R26100 VSS.n4121 VSS.n4120 0.00222973
R26101 VSS.n2514 VSS.n2513 0.00222973
R26102 VSS.n2610 VSS.n1836 0.00222973
R26103 VSS.n2100 VSS.n2097 0.00222973
R26104 VSS.n2771 VSS.n1463 0.00222973
R26105 VSS.n3360 VSS.n3222 0.00222482
R26106 VSS.n3957 VSS.n3936 0.00222482
R26107 VSS.n2275 VSS.n1989 0.00222482
R26108 VSS.n2406 VSS.n1927 0.00222482
R26109 VSS.n3342 VSS.n3229 0.0022027
R26110 VSS.n2250 VSS.n1995 0.0022027
R26111 VSS.n3439 VSS.n3381 0.00220238
R26112 VSS.n3408 VSS.n3407 0.00220238
R26113 VSS.n2304 VSS.n2303 0.00220238
R26114 VSS.n2348 VSS.n1952 0.00220238
R26115 VSS.n3427 VSS.n3388 0.00217619
R26116 VSS.n3422 VSS.n3421 0.00217619
R26117 VSS.n2320 VSS.n2319 0.00217619
R26118 VSS.n2327 VSS.n2326 0.00217619
R26119 VSS.n2783 VSS.n2782 0.00217613
R26120 VSS.n3301 VSS.n3240 0.00215848
R26121 VSS.n3991 VSS.n3920 0.00215848
R26122 VSS.n2214 VSS.n2011 0.00215848
R26123 VSS.n2464 VSS.n1909 0.00215848
R26124 VSS.n3323 VSS.n3233 0.00213636
R26125 VSS.n3970 VSS.n3926 0.00213636
R26126 VSS.n3742 VSS.n3060 0.00213636
R26127 VSS.n3813 VSS.n3032 0.00213636
R26128 VSS.n1707 VSS.n1706 0.00213636
R26129 VSS.n1753 VSS.n1749 0.00213636
R26130 VSS.n2234 VSS.n2003 0.00213636
R26131 VSS.n2419 VSS.n1917 0.00213636
R26132 VSS.n3540 VSS.n3156 0.00211425
R26133 VSS.n3651 VSS.n3103 0.00211425
R26134 VSS.n4088 VSS.n3885 0.00211425
R26135 VSS.n4166 VSS.n3867 0.00211425
R26136 VSS.n2568 VSS.n1859 0.00211425
R26137 VSS.n2670 VSS.n2669 0.00211425
R26138 VSS.n2141 VSS.n2077 0.00211425
R26139 VSS.n1623 VSS.n1570 0.00211425
R26140 VSS.n4037 VSS.n4036 0.00209762
R26141 VSS.n3287 VSS.n3286 0.00209762
R26142 VSS.n2499 VSS.n2498 0.00209762
R26143 VSS.n2200 VSS.n2199 0.00209762
R26144 VSS.n3411 VSS.n3410 0.00209214
R26145 VSS.n3501 VSS.n3180 0.00209214
R26146 VSS.n3124 VSS.n3123 0.00209214
R26147 VSS.n4052 VSS.n3893 0.00209214
R26148 VSS.n4132 VSS.n4128 0.00209214
R26149 VSS.n2345 VSS.n1953 0.00209214
R26150 VSS.n2523 VSS.n2521 0.00209214
R26151 VSS.n2625 VSS.n2624 0.00209214
R26152 VSS.n2119 VSS.n2110 0.00209214
R26153 VSS.n1589 VSS.n1580 0.00209214
R26154 VSS.n4002 VSS.n3912 0.00207143
R26155 VSS.n2451 VSS.n2450 0.00207143
R26156 VSS.n3371 VSS.n3370 0.00207002
R26157 VSS.n3436 VSS.n3382 0.00207002
R26158 VSS.n2288 VSS.n1974 0.00207002
R26159 VSS.n2310 VSS.n1967 0.00207002
R26160 VSS.n4281 VSS.n4280 0.00204791
R26161 VSS.n2362 VSS.n1944 0.00204791
R26162 VSS.n3270 VSS.n3252 0.0020258
R26163 VSS.n4017 VSS.n4016 0.0020258
R26164 VSS.n4027 VSS.n3908 0.0020258
R26165 VSS.n2038 VSS.n2037 0.0020258
R26166 VSS.n2481 VSS.n1900 0.0020258
R26167 VSS.n2483 VSS.n2482 0.0020258
R26168 VSS.n3374 VSS.n3214 0.00201905
R26169 VSS.n2295 VSS.n1973 0.00201905
R26170 VSS.n3496 VSS.n3175 0.00201351
R26171 VSS.n3609 VSS.n3608 0.00201351
R26172 VSS.n4057 VSS.n2969 0.00201351
R26173 VSS.n3873 VSS.n2990 0.00201351
R26174 VSS.n2533 VSS.n2532 0.00201351
R26175 VSS.n2618 VSS.n2617 0.00201351
R26176 VSS.n2112 VSS.n2061 0.00201351
R26177 VSS.n1585 VSS.n1584 0.00201351
R26178 VSS.n3277 VSS.n3274 0.00200369
R26179 VSS.n3248 VSS.n3245 0.00200369
R26180 VSS.n3717 VSS.n3716 0.00200369
R26181 VSS.n3849 VSS.n3848 0.00200369
R26182 VSS.n1670 VSS.n1558 0.00200369
R26183 VSS.n1787 VSS.n1534 0.00200369
R26184 VSS.n2190 VSS.n2024 0.00200369
R26185 VSS.n2020 VSS.n2017 0.00200369
R26186 VSS.n3266 VSS.n3264 0.00200107
R26187 VSS.n3265 VSS.n3192 0.00200107
R26188 VSS.n4033 VSS.n3905 0.00200107
R26189 VSS.n2502 VSS.n2490 0.00200107
R26190 VSS.n2046 VSS.n2045 0.00200107
R26191 VSS.n2169 VSS.n2168 0.00200107
R26192 VSS.n4285 VSS.n4284 0.00199286
R26193 VSS.n2359 VSS.n2358 0.00199286
R26194 VSS.n3999 VSS.n3915 0.00198157
R26195 VSS.n2455 VSS.n2454 0.00198157
R26196 VSS.n1021 VSS.n481 0.00194262
R26197 VSS.n1041 VSS.n473 0.00194262
R26198 VSS.n1058 VSS.n465 0.00194262
R26199 VSS.n1076 VSS.n1067 0.00194262
R26200 VSS.n3438 VSS.n3437 0.00193735
R26201 VSS.n3406 VSS.n3398 0.00193735
R26202 VSS.n2305 VSS.n1970 0.00193735
R26203 VSS.n2347 VSS.n2346 0.00193735
R26204 VSS.n3426 VSS.n3425 0.00191523
R26205 VSS.n3420 VSS.n3392 0.00191523
R26206 VSS.n3267 VSS.n3255 0.00191523
R26207 VSS.n3258 VSS.n3257 0.00191523
R26208 VSS.n4032 VSS.n3907 0.00191523
R26209 VSS.n4186 VSS.n3858 0.00191523
R26210 VSS.n2318 VSS.n1962 0.00191523
R26211 VSS.n2325 VSS.n1963 0.00191523
R26212 VSS.n2503 VSS.n1896 0.00191523
R26213 VSS.n2695 VSS.n1530 0.00191523
R26214 VSS.n2171 VSS.n2033 0.00191523
R26215 VSS.n2170 VSS.n2047 0.00191523
R26216 VSS.n3314 VSS.n3234 0.00191429
R26217 VSS.n3977 VSS.n3925 0.00191429
R26218 VSS.n2228 VSS.n2227 0.00191429
R26219 VSS.n2422 VSS.n1914 0.00191429
R26220 VSS.n672 VSS.n668 0.0019061
R26221 VSS.n3327 VSS.n3326 0.00187101
R26222 VSS.n2239 VSS.n2238 0.00187101
R26223 VSS.n687 VSS.n686 0.00185625
R26224 VSS.n3499 VSS.n3498 0.00185493
R26225 VSS.n3606 VSS.n3121 0.00185493
R26226 VSS.n2117 VSS.n2114 0.00185493
R26227 VSS.n1587 VSS.n1581 0.00185493
R26228 VSS.n3285 VSS.n3247 0.00184889
R26229 VSS.n3969 VSS.n3930 0.00184889
R26230 VSS.n3773 VSS.n3056 0.00184889
R26231 VSS.n3788 VSS.n3042 0.00184889
R26232 VSS.n3475 VSS.n3193 0.00184889
R26233 VSS.n3573 VSS.n3572 0.00184889
R26234 VSS.n3579 VSS.n3143 0.00184889
R26235 VSS.n3682 VSS.n3093 0.00184889
R26236 VSS.n4038 VSS.n3897 0.00184889
R26237 VSS.n4100 VSS.n3880 0.00184889
R26238 VSS.n4115 VSS.n4111 0.00184889
R26239 VSS.n4182 VSS.n4181 0.00184889
R26240 VSS.n1724 VSS.n1723 0.00184889
R26241 VSS.n1733 VSS.n1545 0.00184889
R26242 VSS.n2198 VSS.n2019 0.00184889
R26243 VSS.n2418 VSS.n1920 0.00184889
R26244 VSS.n2497 VSS.n2495 0.00184889
R26245 VSS.n2593 VSS.n2592 0.00184889
R26246 VSS.n2602 VSS.n2601 0.00184889
R26247 VSS.n2692 VSS.n2691 0.00184889
R26248 VSS.n2166 VSS.n2052 0.00184889
R26249 VSS.n2790 VSS.n2789 0.00184889
R26250 VSS.n2778 VSS.n1459 0.00184889
R26251 VSS.n1648 VSS.n1647 0.00184889
R26252 VSS.n3948 VSS.n3937 0.00183571
R26253 VSS.n2397 VSS.n1928 0.00183571
R26254 VSS.n3916 VSS.n3913 0.00182678
R26255 VSS.n2449 VSS.n2444 0.00182678
R26256 VSS.n3346 VSS.n3345 0.00180952
R26257 VSS.n2259 VSS.n1992 0.00180952
R26258 VSS.n3335 VSS.n3226 0.0017973
R26259 VSS.n3952 VSS.n3935 0.0017973
R26260 VSS.n3752 VSS.n3751 0.0017973
R26261 VSS.n3820 VSS.n3027 0.0017973
R26262 VSS.n1695 VSS.n1553 0.0017973
R26263 VSS.n1760 VSS.n1515 0.0017973
R26264 VSS.n2255 VSS.n1994 0.0017973
R26265 VSS.n2401 VSS.n1926 0.0017973
R26266 VSS.n3473 VSS.n3189 0.0017897
R26267 VSS.n3140 VSS.n3139 0.0017897
R26268 VSS.n2164 VSS.n2053 0.0017897
R26269 VSS.n2775 VSS.n2774 0.0017897
R26270 VSS.n3369 VSS.n3218 0.00178256
R26271 VSS.n3376 VSS.n3375 0.00178256
R26272 VSS.n4277 VSS.n2937 0.00178256
R26273 VSS.n2287 VSS.n1977 0.00178256
R26274 VSS.n2294 VSS.n2293 0.00178256
R26275 VSS.n2372 VSS.n2371 0.00178256
R26276 VSS.n4286 VSS.n2934 0.00176044
R26277 VSS.n2360 VSS.n1947 0.00176044
R26278 VSS.n3662 VSS.n3661 0.00175714
R26279 VSS.n1638 VSS.n1637 0.00175714
R26280 VSS.n731 VSS 0.00175595
R26281 VSS.n1003 VSS.n495 0.00175
R26282 VSS.n934 VSS.n756 0.00175
R26283 VSS.n3347 VSS.n3224 0.00173095
R26284 VSS.n3947 VSS.n3946 0.00173095
R26285 VSS.n2261 VSS.n2260 0.00173095
R26286 VSS.n2396 VSS.n2395 0.00173095
R26287 VSS.n3294 VSS.n3293 0.00171622
R26288 VSS.n2207 VSS.n2206 0.00171622
R26289 VSS.n3553 VSS.n3552 0.00171347
R26290 VSS.n2794 VSS.n1456 0.00171347
R26291 VSS.n1100 VSS.n1099 0.00170566
R26292 VSS.n3315 VSS.n3235 0.0016941
R26293 VSS.n3976 VSS.n3975 0.0016941
R26294 VSS.n3998 VSS.n3997 0.0016941
R26295 VSS.n3701 VSS.n3700 0.0016941
R26296 VSS.n4193 VSS.n4192 0.0016941
R26297 VSS.n1664 VSS.n1561 0.0016941
R26298 VSS.n1799 VSS.n1794 0.0016941
R26299 VSS.n2229 VSS.n2005 0.0016941
R26300 VSS.n1918 VSS.n1915 0.0016941
R26301 VSS.n2458 VSS.n2439 0.0016941
R26302 VSS.n3978 VSS.n3923 0.00165238
R26303 VSS.n2431 VSS.n2430 0.00165238
R26304 VSS.n697 VSS.n696 0.00164583
R26305 VSS.n652 VSS.n597 0.00164583
R26306 VSS.n661 VSS.n649 0.00164583
R26307 VSS.n663 VSS.n598 0.00164583
R26308 VSS.n665 VSS.n648 0.00164583
R26309 VSS.n676 VSS.n599 0.00164583
R26310 VSS.n678 VSS.n600 0.00164583
R26311 VSS.n680 VSS.n608 0.00164583
R26312 VSS.n610 VSS.n609 0.00164583
R26313 VSS.n611 VSS.n586 0.00164583
R26314 VSS.n613 VSS.n612 0.00164583
R26315 VSS.n700 VSS.n594 0.00164583
R26316 VSS.n699 VSS.n595 0.00164583
R26317 VSS.n623 VSS.n614 0.00164583
R26318 VSS.n616 VSS.n615 0.00164583
R26319 VSS.n646 VSS.n645 0.00164583
R26320 VSS.n642 VSS.n602 0.00164583
R26321 VSS.n640 VSS.n606 0.00164583
R26322 VSS.n638 VSS.n603 0.00164583
R26323 VSS.n636 VSS.n605 0.00164583
R26324 VSS.n710 VSS.n579 0.00164583
R26325 VSS.n711 VSS.n578 0.00164583
R26326 VSS.n709 VSS.n577 0.00164583
R26327 VSS.n712 VSS.n576 0.00164583
R26328 VSS.n3390 VSS.n3387 0.00162776
R26329 VSS.n3419 VSS.n3417 0.00162776
R26330 VSS.n3949 VSS.n3938 0.00162776
R26331 VSS.n4029 VSS.n3903 0.00162776
R26332 VSS.n2317 VSS.n2316 0.00162776
R26333 VSS.n2324 VSS.n2323 0.00162776
R26334 VSS.n2398 VSS.n1929 0.00162776
R26335 VSS.n2492 VSS.n2491 0.00162776
R26336 VSS.n3313 VSS.n3312 0.00162619
R26337 VSS.n2226 VSS.n2225 0.00162619
R26338 VSS.n3344 VSS.n3227 0.00160565
R26339 VSS.n2258 VSS.n1993 0.00160565
R26340 VSS.n3478 VSS.n3187 0.00158354
R26341 VSS.n3600 VSS.n3599 0.00158354
R26342 VSS.n4045 VSS.n3896 0.00158354
R26343 VSS.n4119 VSS.n4118 0.00158354
R26344 VSS.n2516 VSS.n2515 0.00158354
R26345 VSS.n1844 VSS.n1843 0.00158354
R26346 VSS.n2101 VSS.n2099 0.00158354
R26347 VSS.n2770 VSS.n1462 0.00158354
R26348 VSS.n3284 VSS.n3283 0.00156143
R26349 VSS.n4008 VSS.n4007 0.00156143
R26350 VSS.n3770 VSS.n3769 0.00156143
R26351 VSS.n3792 VSS.n3791 0.00156143
R26352 VSS.n3557 VSS.n3556 0.00156143
R26353 VSS.n3660 VSS.n3659 0.00156143
R26354 VSS.n4097 VSS.n4096 0.00156143
R26355 VSS.n4175 VSS.n4174 0.00156143
R26356 VSS.n1715 VSS.n1548 0.00156143
R26357 VSS.n1740 VSS.n1543 0.00156143
R26358 VSS.n2197 VSS.n2196 0.00156143
R26359 VSS.n2448 VSS.n2447 0.00156143
R26360 VSS.n2574 VSS.n2573 0.00156143
R26361 VSS.n2679 VSS.n2678 0.00156143
R26362 VSS.n2796 VSS.n1452 0.00156143
R26363 VSS.n1639 VSS.n1565 0.00156143
R26364 VSS.n3380 VSS.n3379 0.00154762
R26365 VSS.n3402 VSS.n2935 0.00154762
R26366 VSS.n2296 VSS.n1971 0.00154762
R26367 VSS.n2357 VSS.n1948 0.00154762
R26368 VSS.n3348 VSS.n3225 0.00153931
R26369 VSS.n3945 VSS.n3939 0.00153931
R26370 VSS.n2262 VSS.n1991 0.00153931
R26371 VSS.n2394 VSS.n1931 0.00153931
R26372 VSS.n571 VSS.n570 0.00153774
R26373 VSS.n567 VSS.n524 0.00153774
R26374 VSS.n565 VSS.n530 0.00153774
R26375 VSS.n563 VSS.n525 0.00153774
R26376 VSS.n561 VSS.n529 0.00153774
R26377 VSS.n559 VSS.n527 0.00153774
R26378 VSS.n957 VSS.n522 0.00153774
R26379 VSS.n956 VSS.n518 0.00153774
R26380 VSS.n961 VSS.n958 0.00153774
R26381 VSS.n960 VSS.n517 0.00153774
R26382 VSS.n963 VSS.n515 0.00153774
R26383 VSS.n965 VSS.n964 0.00153774
R26384 VSS.n967 VSS.n501 0.00153774
R26385 VSS.n969 VSS.n502 0.00153774
R26386 VSS.n504 VSS.n503 0.00153774
R26387 VSS.n1000 VSS.n999 0.00153774
R26388 VSS.n996 VSS.n496 0.00153774
R26389 VSS.n994 VSS.n500 0.00153774
R26390 VSS.n992 VSS.n497 0.00153774
R26391 VSS.n990 VSS.n499 0.00153774
R26392 VSS.n1178 VSS.n1157 0.00152655
R26393 VSS.n836 VSS.n760 0.00152255
R26394 VSS.n3378 VSS.n3377 0.00149509
R26395 VSS.n3658 VSS.n3657 0.00149509
R26396 VSS.n2297 VSS.n1972 0.00149509
R26397 VSS.n1625 VSS.n1566 0.00149509
R26398 VSS.n4287 VSS.n2933 0.00147297
R26399 VSS.n3980 VSS.n3979 0.00147297
R26400 VSS.n2356 VSS.n2355 0.00147297
R26401 VSS.n2429 VSS.n1912 0.00147297
R26402 VSS.n3281 VSS.n3249 0.00146905
R26403 VSS.n4010 VSS.n4009 0.00146905
R26404 VSS.n2194 VSS.n2021 0.00146905
R26405 VSS.n2446 VSS.n2445 0.00146905
R26406 VSS.n3311 VSS.n3236 0.00145086
R26407 VSS.n2224 VSS.n2007 0.00145086
R26408 VSS.n3316 VSS.n3236 0.00140663
R26409 VSS.n3979 VSS.n3924 0.00140663
R26410 VSS.n3713 VSS.n3712 0.00140663
R26411 VSS.n3834 VSS.n3016 0.00140663
R26412 VSS.n1677 VSS.n1556 0.00140663
R26413 VSS.n1780 VSS.n1535 0.00140663
R26414 VSS.n2230 VSS.n2007 0.00140663
R26415 VSS.n2429 VSS.n2428 0.00140663
R26416 VSS.n3415 VSS.n3393 0.00139048
R26417 VSS.n2322 VSS.n2321 0.00139048
R26418 VSS.n3378 VSS.n3212 0.00138452
R26419 VSS.n3401 VSS.n2933 0.00138452
R26420 VSS.n2298 VSS.n2297 0.00138452
R26421 VSS.n2356 VSS.n1949 0.00138452
R26422 VSS.n3273 VSS.n3272 0.00136429
R26423 VSS.n3435 VSS.n3381 0.00136429
R26424 VSS.n3429 VSS.n3428 0.00136429
R26425 VSS.n2036 VSS.n2035 0.00136429
R26426 VSS.n2303 VSS.n2302 0.00136429
R26427 VSS.n2314 VSS.n1964 0.00136429
R26428 VSS.n3349 VSS.n3348 0.00134029
R26429 VSS.n3950 VSS.n3939 0.00134029
R26430 VSS.n2257 VSS.n1991 0.00134029
R26431 VSS.n2399 VSS.n1931 0.00134029
R26432 VSS.n3409 VSS.n3408 0.00133809
R26433 VSS.n4019 VSS.n4018 0.00133809
R26434 VSS.n2344 VSS.n1952 0.00133809
R26435 VSS.n2480 VSS.n1899 0.00133809
R26436 VSS.n3283 VSS.n3282 0.00131818
R26437 VSS.n4008 VSS.n3911 0.00131818
R26438 VSS.n3556 VSS.n3555 0.00131818
R26439 VSS.n2196 VSS.n2195 0.00131818
R26440 VSS.n2447 VSS.n1902 0.00131818
R26441 VSS.n2796 VSS.n2795 0.00131818
R26442 VSS.n4059 VSS.n3892 0.00129607
R26443 VSS.n4081 VSS.n3887 0.00129607
R26444 VSS.n4136 VSS.n4135 0.00129607
R26445 VSS.n4159 VSS.n3868 0.00129607
R26446 VSS.n2538 VSS.n2537 0.00129607
R26447 VSS.n2562 VSS.n2561 0.00129607
R26448 VSS.n2621 VSS.n2620 0.00129607
R26449 VSS.n2654 VSS.n2651 0.00129607
R26450 VSS.n1099 VSS.n454 0.00129432
R26451 VSS.n3296 VSS.n3295 0.00128571
R26452 VSS.n3995 VSS.n3917 0.00128571
R26453 VSS.n2209 VSS.n2208 0.00128571
R26454 VSS.n2457 VSS.n2438 0.00128571
R26455 VSS.n3349 VSS.n3227 0.00125184
R26456 VSS.n3417 VSS.n3416 0.00125184
R26457 VSS.n3950 VSS.n3949 0.00125184
R26458 VSS.n3748 VSS.n3069 0.00125184
R26459 VSS.n3817 VSS.n3816 0.00125184
R26460 VSS.n1699 VSS.n1698 0.00125184
R26461 VSS.n1757 VSS.n1756 0.00125184
R26462 VSS.n2258 VSS.n2257 0.00125184
R26463 VSS.n2323 VSS.n1955 0.00125184
R26464 VSS.n2399 VSS.n2398 0.00125184
R26465 VSS.n1003 VSS.n1002 0.00124998
R26466 VSS.n3274 VSS.n3252 0.00122973
R26467 VSS.n3437 VSS.n3436 0.00122973
R26468 VSS.n3430 VSS.n3387 0.00122973
R26469 VSS.n2037 VSS.n2024 0.00122973
R26470 VSS.n1970 VSS.n1967 0.00122973
R26471 VSS.n2316 VSS.n2315 0.00122973
R26472 VSS.n3410 VSS.n3398 0.00120762
R26473 VSS.n4017 VSS.n3908 0.00120762
R26474 VSS.n2346 VSS.n2345 0.00120762
R26475 VSS.n2482 VSS.n2481 0.00120762
R26476 VSS.n3364 VSS.n3363 0.00120714
R26477 VSS.n4278 VSS.n2938 0.00120714
R26478 VSS.n2268 VSS.n1976 0.00120714
R26479 VSS.n2370 VSS.n2369 0.00120714
R26480 VSS.n3316 VSS.n3315 0.0011855
R26481 VSS.n3976 VSS.n3924 0.0011855
R26482 VSS.n2230 VSS.n2229 0.0011855
R26483 VSS.n2428 VSS.n1915 0.0011855
R26484 VSS.n672 VSS.n670 0.00116947
R26485 VSS.n3294 VSS.n3243 0.00116339
R26486 VSS.n3997 VSS.n3996 0.00116339
R26487 VSS.n2207 VSS.n2015 0.00116339
R26488 VSS.n2459 VSS.n2458 0.00116339
R26489 VSS.n3490 VSS.n3185 0.00114865
R26490 VSS.n3594 VSS.n3590 0.00114865
R26491 VSS.n4049 VSS.n4048 0.00114865
R26492 VSS.n4123 VSS.n2988 0.00114865
R26493 VSS.n2526 VSS.n1883 0.00114865
R26494 VSS.n2613 VSS.n2612 0.00114865
R26495 VSS.n2104 VSS.n2059 0.00114865
R26496 VSS.n2767 VSS.n1465 0.00114865
R26497 VSS.n3964 VSS.n3929 0.00112857
R26498 VSS.n2413 VSS.n1919 0.00112857
R26499 VSS.n4287 VSS.n4286 0.00111916
R26500 VSS.n2355 VSS.n1947 0.00111916
R26501 VSS.n3329 VSS.n3232 0.00110238
R26502 VSS.n2237 VSS.n2000 0.00110238
R26503 VSS.n3220 VSS.n3218 0.00109705
R26504 VSS.n3377 VSS.n3376 0.00109705
R26505 VSS.n4277 VSS.n4276 0.00109705
R26506 VSS.n3750 VSS.n3068 0.00109705
R26507 VSS.n3822 VSS.n3821 0.00109705
R26508 VSS.n3657 VSS.n3654 0.00109705
R26509 VSS.n1694 VSS.n1693 0.00109705
R26510 VSS.n1762 VSS.n1761 0.00109705
R26511 VSS.n2269 VSS.n1977 0.00109705
R26512 VSS.n2294 VSS.n1972 0.00109705
R26513 VSS.n2371 VSS.n1945 0.00109705
R26514 VSS.n1625 VSS.n1567 0.00109705
R26515 VSS.n4077 VSS.n4076 0.00105283
R26516 VSS.n4155 VSS.n4154 0.00105283
R26517 VSS.n4189 VSS.n3858 0.00105283
R26518 VSS.n2542 VSS.n1864 0.00105283
R26519 VSS.n2656 VSS.n2649 0.00105283
R26520 VSS.n1802 VSS.n1530 0.00105283
R26521 VSS.n3389 VSS.n2928 0.00104054
R26522 VSS.n3054 VSS.n3053 0.00104054
R26523 VSS.n1721 VSS.n1506 0.00104054
R26524 VSS.n2331 VSS.n1960 0.00104054
R26525 VSS.n3285 VSS.n3284 0.00103071
R26526 VSS.n3932 VSS.n3930 0.00103071
R26527 VSS.n4007 VSS.n3913 0.00103071
R26528 VSS.n3262 VSS.n3255 0.00103071
R26529 VSS.n3475 VSS.n3474 0.00103071
R26530 VSS.n3143 VSS.n3142 0.00103071
R26531 VSS.n4022 VSS.n3907 0.00103071
R26532 VSS.n4062 VSS.n4061 0.00103071
R26533 VSS.n4142 VSS.n4141 0.00103071
R26534 VSS.n2198 VSS.n2197 0.00103071
R26535 VSS.n1923 VSS.n1920 0.00103071
R26536 VSS.n2449 VSS.n2448 0.00103071
R26537 VSS.n2488 VSS.n1896 0.00103071
R26538 VSS.n1877 VSS.n1871 0.00103071
R26539 VSS.n2639 VSS.n2638 0.00103071
R26540 VSS.n2043 VSS.n2033 0.00103071
R26541 VSS.n2166 VSS.n2165 0.00103071
R26542 VSS.n1460 VSS.n1459 0.00103071
R26543 VSS.n1255 VSS.n1254 0.00102242
R26544 VSS.n3328 VSS.n3327 0.0010086
R26545 VSS.n2238 VSS.n2001 0.0010086
R26546 VSS.n1095 VSS.n1094 0.00100303
R26547 VSS.n454 VSS.n451 0.001
R26548 VSS.n1114 VSS.n1113 0.001
R26549 VSS.n955 VSS.n493 0.001
R26550 VSS.n959 VSS.n494 0.001
R26551 VSS.n495 VSS.n494 0.001
R26552 VSS.n959 VSS.n493 0.001
R26553 VSS.n1130 VSS.n1114 0.001
R26554 VSS.n1100 VSS.n451 0.001
R26555 VSS.n3426 VSS.n3390 0.000964373
R26556 VSS.n3420 VSS.n3419 0.000964373
R26557 VSS.n3257 VSS.n3256 0.000964373
R26558 VSS.n3688 VSS.n3687 0.000964373
R26559 VSS.n4029 VSS.n3904 0.000964373
R26560 VSS.n2318 VSS.n2317 0.000964373
R26561 VSS.n2325 VSS.n2324 0.000964373
R26562 VSS.n2491 VSS.n1897 0.000964373
R26563 VSS.n2048 VSS.n2047 0.000964373
R26564 VSS.n1644 VSS.n1563 0.000964373
R26565 VSS.n3730 VSS.n3729 0.00094226
R26566 VSS.n3836 VSS.n3833 0.00094226
R26567 VSS.n1682 VSS.n1681 0.00094226
R26568 VSS.n1776 VSS.n1775 0.00094226
R26569 VSS.n3186 VSS.n3181 0.000932432
R26570 VSS.n3591 VSS.n3122 0.000932432
R26571 VSS.n4053 VSS.n2968 0.000932432
R26572 VSS.n4129 VSS.n2989 0.000932432
R26573 VSS.n2522 VSS.n1884 0.000932432
R26574 VSS.n2627 VSS.n2626 0.000932432
R26575 VSS.n2115 VSS.n2060 0.000932432
R26576 VSS.n2762 VSS.n1469 0.000932432
R26577 VSS.n3267 VSS.n3254 0.000898034
R26578 VSS.n3999 VSS.n3998 0.000898034
R26579 VSS.n2171 VSS.n2032 0.000898034
R26580 VSS.n2455 VSS.n2439 0.000898034
R26581 VSS.n3293 VSS.n3245 0.000875921
R26582 VSS.n2206 VSS.n2017 0.000875921
R26583 VSS.n1022 VSS.n1021 0.000860656
R26584 VSS.n1042 VSS.n1041 0.000860656
R26585 VSS.n1059 VSS.n1058 0.000860656
R26586 VSS.n1076 VSS.n455 0.000860656
R26587 VSS.n1098 VSS.n1097 0.000860656
R26588 VSS.n4032 VSS.n3906 0.000853808
R26589 VSS.n2503 VSS.n1895 0.000853808
R26590 VSS.n725 VSS.n724 0.000834919
R26591 VSS.n721 VSS.n718 0.000834919
R26592 VSS.n3669 VSS.n3668 0.000831695
R26593 VSS.n1631 VSS.n1630 0.000831695
R26594 VSS.n3666 VSS.n3665 0.000814286
R26595 VSS.n1634 VSS.n1633 0.000814286
R26596 VSS.n3370 VSS.n3369 0.000809582
R26597 VSS.n4280 VSS.n2937 0.000809582
R26598 VSS.n2288 VSS.n2287 0.000809582
R26599 VSS.n2372 VSS.n1944 0.000809582
R26600 VSS.n3764 VSS.n3763 0.000787469
R26601 VSS.n3797 VSS.n3796 0.000787469
R26602 VSS.n3501 VSS.n3500 0.000787469
R26603 VSS.n3605 VSS.n3123 0.000787469
R26604 VSS.n1711 VSS.n1710 0.000787469
R26605 VSS.n1745 VSS.n1744 0.000787469
R26606 VSS.n2119 VSS.n2118 0.000787469
R26607 VSS.n1589 VSS.n1588 0.000787469
R26608 VSS.n3653 VSS.n3104 0.000765356
R26609 VSS.n4047 VSS.n3894 0.000765356
R26610 VSS.n4092 VSS.n3884 0.000765356
R26611 VSS.n4125 VSS.n4124 0.000765356
R26612 VSS.n4171 VSS.n4170 0.000765356
R26613 VSS.n2519 VSS.n1885 0.000765356
R26614 VSS.n2577 VSS.n1860 0.000765356
R26615 VSS.n2615 VSS.n2614 0.000765356
R26616 VSS.n2674 VSS.n2673 0.000765356
R26617 VSS.n1632 VSS.n1568 0.000765356
R26618 VSS.n3970 VSS.n3969 0.000743243
R26619 VSS.n2419 VSS.n2418 0.000743243
R26620 VSS.n3326 VSS.n3323 0.00072113
R26621 VSS.n2239 VSS.n2003 0.00072113
R26622 VSS.n3292 VSS.n3199 0.000716216
R26623 VSS.n3914 VSS.n2958 0.000716216
R26624 VSS.n3719 VSS.n3080 0.000716216
R26625 VSS.n3852 VSS.n3851 0.000716216
R26626 VSS.n1668 VSS.n1492 0.000716216
R26627 VSS.n1790 VSS.n1521 0.000716216
R26628 VSS.n2205 VSS.n2014 0.000716216
R26629 VSS.n2442 VSS.n2441 0.000716216
R26630 VSS.n3337 VSS.n3229 0.000676904
R26631 VSS.n2250 VSS.n2249 0.000676904
R26632 VSS.n734 VSS.n713 0.00066746
R26633 VSS.n733 VSS.n714 0.00066746
R26634 VSS.n725 VSS.n714 0.00066746
R26635 VSS.n724 VSS.n717 0.00066746
R26636 VSS.n730 VSS.n729 0.00066746
R26637 VSS.n729 VSS.n718 0.00066746
R26638 VSS.n721 VSS.n516 0.00066746
R26639 VSS.n3958 VSS.n3957 0.000654791
R26640 VSS.n3707 VSS.n3706 0.000654791
R26641 VSS.n3855 VSS.n3854 0.000654791
R26642 VSS.n1666 VSS.n1559 0.000654791
R26643 VSS.n1788 VSS.n1533 0.000654791
R26644 VSS.n2407 VSS.n2406 0.000654791
R26645 VSS.n4269 VSS.n2945 0.000588452
R26646 VSS.n2387 VSS.n1933 0.000588452
R26647 VSS.n962 VSS.n513 0.00058373
R26648 VSS.n3357 VSS.n3356 0.000566339
R26649 VSS.n2276 VSS.n1988 0.000566339
R26650 VSS.n3307 VSS.n3306 0.000522113
R26651 VSS.n3094 VSS.n3087 0.000522113
R26652 VSS.n1657 VSS.n1562 0.000522113
R26653 VSS.n2220 VSS.n2219 0.000522113
R26654 VDD.n74 VDD.n71 17.001
R26655 VDD.n305 VDD.n304 17.0005
R26656 VDD.n299 VDD.n294 17.0005
R26657 VDD.n310 VDD.n284 17.0005
R26658 VDD.n2045 VDD.n2041 17.0005
R26659 VDD.n2037 VDD.n2036 17.0005
R26660 VDD.n2028 VDD.n2019 17.0005
R26661 VDD.n1937 VDD.n565 12.5814
R26662 VDD.n1938 VDD 12.1116
R26663 VDD.n302 VDD.n301 10.9321
R26664 VDD.n302 VDD.n293 10.9321
R26665 VDD.n2039 VDD.n2038 10.9321
R26666 VDD.n2039 VDD.n2029 10.9321
R26667 VDD.n579 VDD 9.14886
R26668 VDD.n561 VDD.n560 9.10654
R26669 VDD.n556 VDD.n555 9.10333
R26670 VDD.n560 VDD.n555 9.10238
R26671 VDD.n442 VDD.n441 9.07498
R26672 VDD.n523 VDD.n522 9.07375
R26673 VDD.n85 VDD.n84 9.05588
R26674 VDD.n569 VDD.n567 9.04906
R26675 VDD.n572 VDD.n566 9.049
R26676 VDD.n579 VDD.n578 9.03124
R26677 VDD.n578 VDD.n577 9.03024
R26678 VDD.n571 VDD.n570 9.0005
R26679 VDD.n573 VDD.n568 9.0005
R26680 VDD.n572 VDD.n571 9.0005
R26681 VDD.n574 VDD.n573 9.0005
R26682 VDD.n575 VDD.n567 9.0005
R26683 VDD.n576 VDD.n575 9.0005
R26684 VDD.n581 VDD.n580 9.0005
R26685 VDD.n559 VDD.n558 9.0005
R26686 VDD.n554 VDD.n553 9.0005
R26687 VDD.n563 VDD.n562 9.0005
R26688 VDD.n558 VDD.n557 9.0005
R26689 VDD.n553 VDD.n552 9.0005
R26690 VDD.n564 VDD.n563 9.0005
R26691 VDD.n552 VDD.n551 9.0005
R26692 VDD.n565 VDD.n564 9.0005
R26693 VDD.n542 VDD.n541 9.0005
R26694 VDD.n543 VDD.n403 9.0005
R26695 VDD.n490 VDD.n401 9.0005
R26696 VDD.n547 VDD.n400 9.0005
R26697 VDD.n548 VDD.n399 9.0005
R26698 VDD.n549 VDD.n398 9.0005
R26699 VDD.n483 VDD.n397 9.0005
R26700 VDD.n482 VDD.n481 9.0005
R26701 VDD.n413 VDD.n412 9.0005
R26702 VDD.n477 VDD.n476 9.0005
R26703 VDD.n416 VDD.n415 9.0005
R26704 VDD.n469 VDD.n468 9.0005
R26705 VDD.n422 VDD.n421 9.0005
R26706 VDD.n464 VDD.n463 9.0005
R26707 VDD.n425 VDD.n424 9.0005
R26708 VDD.n405 VDD.n404 9.0005
R26709 VDD.n541 VDD.n540 9.0005
R26710 VDD.n406 VDD.n403 9.0005
R26711 VDD.n491 VDD.n490 9.0005
R26712 VDD.n489 VDD.n400 9.0005
R26713 VDD.n488 VDD.n399 9.0005
R26714 VDD.n409 VDD.n398 9.0005
R26715 VDD.n484 VDD.n483 9.0005
R26716 VDD.n482 VDD.n411 9.0005
R26717 VDD.n418 VDD.n412 9.0005
R26718 VDD.n476 VDD.n475 9.0005
R26719 VDD.n417 VDD.n416 9.0005
R26720 VDD.n470 VDD.n469 9.0005
R26721 VDD.n421 VDD.n420 9.0005
R26722 VDD.n463 VDD.n462 9.0005
R26723 VDD.n426 VDD.n425 9.0005
R26724 VDD.n407 VDD.n405 9.0005
R26725 VDD.n505 VDD.n504 9.0005
R26726 VDD.n520 VDD.n502 9.0005
R26727 VDD.n519 VDD.n501 9.0005
R26728 VDD.n518 VDD.n500 9.0005
R26729 VDD.n508 VDD.n507 9.0005
R26730 VDD.n514 VDD.n497 9.0005
R26731 VDD.n513 VDD.n496 9.0005
R26732 VDD.n512 VDD.n495 9.0005
R26733 VDD.n504 VDD.n503 9.0005
R26734 VDD.n528 VDD.n502 9.0005
R26735 VDD.n529 VDD.n501 9.0005
R26736 VDD.n530 VDD.n500 9.0005
R26737 VDD.n507 VDD.n498 9.0005
R26738 VDD.n534 VDD.n497 9.0005
R26739 VDD.n535 VDD.n496 9.0005
R26740 VDD.n536 VDD.n495 9.0005
R26741 VDD.n524 VDD.n523 9.0005
R26742 VDD.n525 VDD.n524 9.0005
R26743 VDD.n460 VDD.n426 9.0005
R26744 VDD.n462 VDD.n461 9.0005
R26745 VDD.n420 VDD.n419 9.0005
R26746 VDD.n471 VDD.n470 9.0005
R26747 VDD.n472 VDD.n417 9.0005
R26748 VDD.n475 VDD.n474 9.0005
R26749 VDD.n473 VDD.n418 9.0005
R26750 VDD.n411 VDD.n410 9.0005
R26751 VDD.n485 VDD.n484 9.0005
R26752 VDD.n486 VDD.n409 9.0005
R26753 VDD.n488 VDD.n487 9.0005
R26754 VDD.n489 VDD.n408 9.0005
R26755 VDD.n492 VDD.n491 9.0005
R26756 VDD.n493 VDD.n406 9.0005
R26757 VDD.n540 VDD.n539 9.0005
R26758 VDD.n538 VDD.n407 9.0005
R26759 VDD.n537 VDD.n536 9.0005
R26760 VDD.n535 VDD.n494 9.0005
R26761 VDD.n534 VDD.n533 9.0005
R26762 VDD.n532 VDD.n498 9.0005
R26763 VDD.n531 VDD.n530 9.0005
R26764 VDD.n529 VDD.n499 9.0005
R26765 VDD.n528 VDD.n527 9.0005
R26766 VDD.n526 VDD.n503 9.0005
R26767 VDD.n440 VDD.n439 9.0005
R26768 VDD.n436 VDD.n435 9.0005
R26769 VDD.n447 VDD.n446 9.0005
R26770 VDD.n448 VDD.n434 9.0005
R26771 VDD.n450 VDD.n449 9.0005
R26772 VDD.n428 VDD.n427 9.0005
R26773 VDD.n459 VDD.n458 9.0005
R26774 VDD.n429 VDD.n428 9.0005
R26775 VDD.n451 VDD.n450 9.0005
R26776 VDD.n434 VDD.n433 9.0005
R26777 VDD.n446 VDD.n445 9.0005
R26778 VDD.n437 VDD.n436 9.0005
R26779 VDD.n441 VDD.n440 9.0005
R26780 VDD.n458 VDD.n457 9.0005
R26781 VDD.n430 VDD.n429 9.0005
R26782 VDD.n452 VDD.n451 9.0005
R26783 VDD.n433 VDD.n432 9.0005
R26784 VDD.n445 VDD.n444 9.0005
R26785 VDD.n438 VDD.n437 9.0005
R26786 VDD.n457 VDD.n456 9.0005
R26787 VDD.n454 VDD.n430 9.0005
R26788 VDD.n453 VDD.n452 9.0005
R26789 VDD.n432 VDD.n431 9.0005
R26790 VDD.n444 VDD.n443 9.0005
R26791 VDD.n456 VDD.n455 9.0005
R26792 VDD.n542 VDD.n402 9.0005
R26793 VDD.n544 VDD.n543 9.0005
R26794 VDD.n545 VDD.n401 9.0005
R26795 VDD.n547 VDD.n546 9.0005
R26796 VDD.n548 VDD.n396 9.0005
R26797 VDD.n550 VDD.n549 9.0005
R26798 VDD.n397 VDD.n395 9.0005
R26799 VDD.n481 VDD.n480 9.0005
R26800 VDD.n479 VDD.n413 9.0005
R26801 VDD.n478 VDD.n477 9.0005
R26802 VDD.n415 VDD.n414 9.0005
R26803 VDD.n468 VDD.n467 9.0005
R26804 VDD.n466 VDD.n422 9.0005
R26805 VDD.n465 VDD.n464 9.0005
R26806 VDD.n424 VDD.n423 9.0005
R26807 VDD.n510 VDD.n404 9.0005
R26808 VDD.n521 VDD.n520 9.0005
R26809 VDD.n519 VDD.n506 9.0005
R26810 VDD.n518 VDD.n517 9.0005
R26811 VDD.n516 VDD.n508 9.0005
R26812 VDD.n515 VDD.n514 9.0005
R26813 VDD.n513 VDD.n509 9.0005
R26814 VDD.n512 VDD.n511 9.0005
R26815 VDD.n303 VDD.n302 9.0005
R26816 VDD.n313 VDD.n312 9.0005
R26817 VDD.n314 VDD.n278 9.0005
R26818 VDD.n316 VDD.n315 9.0005
R26819 VDD.n318 VDD.n277 9.0005
R26820 VDD.n320 VDD.n319 9.0005
R26821 VDD.n321 VDD.n276 9.0005
R26822 VDD.n323 VDD.n322 9.0005
R26823 VDD.n325 VDD.n275 9.0005
R26824 VDD.n327 VDD.n326 9.0005
R26825 VDD.n328 VDD.n274 9.0005
R26826 VDD.n330 VDD.n329 9.0005
R26827 VDD.n332 VDD.n273 9.0005
R26828 VDD.n334 VDD.n333 9.0005
R26829 VDD.n335 VDD.n272 9.0005
R26830 VDD.n337 VDD.n336 9.0005
R26831 VDD.n339 VDD.n271 9.0005
R26832 VDD.n341 VDD.n340 9.0005
R26833 VDD.n342 VDD.n270 9.0005
R26834 VDD.n344 VDD.n343 9.0005
R26835 VDD.n346 VDD.n269 9.0005
R26836 VDD.n348 VDD.n347 9.0005
R26837 VDD.n349 VDD.n268 9.0005
R26838 VDD.n351 VDD.n350 9.0005
R26839 VDD.n353 VDD.n267 9.0005
R26840 VDD.n355 VDD.n354 9.0005
R26841 VDD.n356 VDD.n266 9.0005
R26842 VDD.n358 VDD.n357 9.0005
R26843 VDD.n360 VDD.n265 9.0005
R26844 VDD.n362 VDD.n361 9.0005
R26845 VDD.n363 VDD.n264 9.0005
R26846 VDD.n365 VDD.n364 9.0005
R26847 VDD.n367 VDD.n263 9.0005
R26848 VDD.n369 VDD.n368 9.0005
R26849 VDD.n370 VDD.n262 9.0005
R26850 VDD.n372 VDD.n371 9.0005
R26851 VDD.n374 VDD.n261 9.0005
R26852 VDD.n376 VDD.n375 9.0005
R26853 VDD.n377 VDD.n260 9.0005
R26854 VDD.n379 VDD.n378 9.0005
R26855 VDD.n381 VDD.n259 9.0005
R26856 VDD.n383 VDD.n382 9.0005
R26857 VDD.n384 VDD.n258 9.0005
R26858 VDD.n386 VDD.n385 9.0005
R26859 VDD.n388 VDD.n257 9.0005
R26860 VDD.n390 VDD.n389 9.0005
R26861 VDD.n391 VDD.n251 9.0005
R26862 VDD.n393 VDD.n392 9.0005
R26863 VDD.n312 VDD.n194 9.0005
R26864 VDD.n278 VDD.n195 9.0005
R26865 VDD.n316 VDD.n196 9.0005
R26866 VDD.n318 VDD.n317 9.0005
R26867 VDD.n319 VDD.n199 9.0005
R26868 VDD.n276 VDD.n200 9.0005
R26869 VDD.n323 VDD.n201 9.0005
R26870 VDD.n325 VDD.n324 9.0005
R26871 VDD.n326 VDD.n204 9.0005
R26872 VDD.n274 VDD.n205 9.0005
R26873 VDD.n330 VDD.n206 9.0005
R26874 VDD.n332 VDD.n331 9.0005
R26875 VDD.n333 VDD.n209 9.0005
R26876 VDD.n272 VDD.n210 9.0005
R26877 VDD.n337 VDD.n211 9.0005
R26878 VDD.n339 VDD.n338 9.0005
R26879 VDD.n340 VDD.n214 9.0005
R26880 VDD.n270 VDD.n215 9.0005
R26881 VDD.n344 VDD.n216 9.0005
R26882 VDD.n346 VDD.n345 9.0005
R26883 VDD.n347 VDD.n219 9.0005
R26884 VDD.n268 VDD.n220 9.0005
R26885 VDD.n351 VDD.n221 9.0005
R26886 VDD.n353 VDD.n352 9.0005
R26887 VDD.n354 VDD.n224 9.0005
R26888 VDD.n266 VDD.n225 9.0005
R26889 VDD.n358 VDD.n226 9.0005
R26890 VDD.n360 VDD.n359 9.0005
R26891 VDD.n361 VDD.n229 9.0005
R26892 VDD.n264 VDD.n230 9.0005
R26893 VDD.n365 VDD.n231 9.0005
R26894 VDD.n367 VDD.n366 9.0005
R26895 VDD.n368 VDD.n234 9.0005
R26896 VDD.n262 VDD.n235 9.0005
R26897 VDD.n372 VDD.n236 9.0005
R26898 VDD.n374 VDD.n373 9.0005
R26899 VDD.n375 VDD.n239 9.0005
R26900 VDD.n260 VDD.n240 9.0005
R26901 VDD.n379 VDD.n241 9.0005
R26902 VDD.n381 VDD.n380 9.0005
R26903 VDD.n382 VDD.n244 9.0005
R26904 VDD.n258 VDD.n245 9.0005
R26905 VDD.n386 VDD.n246 9.0005
R26906 VDD.n388 VDD.n387 9.0005
R26907 VDD.n389 VDD.n249 9.0005
R26908 VDD.n251 VDD.n250 9.0005
R26909 VDD.n394 VDD.n393 9.0005
R26910 VDD.n2009 VDD.n194 9.0005
R26911 VDD.n2008 VDD.n195 9.0005
R26912 VDD.n2007 VDD.n196 9.0005
R26913 VDD.n317 VDD.n197 9.0005
R26914 VDD.n2003 VDD.n199 9.0005
R26915 VDD.n2002 VDD.n200 9.0005
R26916 VDD.n2001 VDD.n201 9.0005
R26917 VDD.n324 VDD.n202 9.0005
R26918 VDD.n1997 VDD.n204 9.0005
R26919 VDD.n1996 VDD.n205 9.0005
R26920 VDD.n1995 VDD.n206 9.0005
R26921 VDD.n331 VDD.n207 9.0005
R26922 VDD.n1991 VDD.n209 9.0005
R26923 VDD.n1990 VDD.n210 9.0005
R26924 VDD.n1989 VDD.n211 9.0005
R26925 VDD.n338 VDD.n212 9.0005
R26926 VDD.n1985 VDD.n214 9.0005
R26927 VDD.n1984 VDD.n215 9.0005
R26928 VDD.n1983 VDD.n216 9.0005
R26929 VDD.n345 VDD.n217 9.0005
R26930 VDD.n1979 VDD.n219 9.0005
R26931 VDD.n1978 VDD.n220 9.0005
R26932 VDD.n1977 VDD.n221 9.0005
R26933 VDD.n352 VDD.n222 9.0005
R26934 VDD.n1973 VDD.n224 9.0005
R26935 VDD.n1972 VDD.n225 9.0005
R26936 VDD.n1971 VDD.n226 9.0005
R26937 VDD.n359 VDD.n227 9.0005
R26938 VDD.n1967 VDD.n229 9.0005
R26939 VDD.n1966 VDD.n230 9.0005
R26940 VDD.n1965 VDD.n231 9.0005
R26941 VDD.n366 VDD.n232 9.0005
R26942 VDD.n1961 VDD.n234 9.0005
R26943 VDD.n1960 VDD.n235 9.0005
R26944 VDD.n1959 VDD.n236 9.0005
R26945 VDD.n373 VDD.n237 9.0005
R26946 VDD.n1955 VDD.n239 9.0005
R26947 VDD.n1954 VDD.n240 9.0005
R26948 VDD.n1953 VDD.n241 9.0005
R26949 VDD.n380 VDD.n242 9.0005
R26950 VDD.n1949 VDD.n244 9.0005
R26951 VDD.n1948 VDD.n245 9.0005
R26952 VDD.n1947 VDD.n246 9.0005
R26953 VDD.n387 VDD.n247 9.0005
R26954 VDD.n1943 VDD.n249 9.0005
R26955 VDD.n1942 VDD.n250 9.0005
R26956 VDD.n1941 VDD.n394 9.0005
R26957 VDD.n49 VDD.n48 9.0005
R26958 VDD.n128 VDD.n127 9.0005
R26959 VDD.n46 VDD.n45 9.0005
R26960 VDD.n133 VDD.n132 9.0005
R26961 VDD.n41 VDD.n40 9.0005
R26962 VDD.n140 VDD.n139 9.0005
R26963 VDD.n38 VDD.n37 9.0005
R26964 VDD.n145 VDD.n144 9.0005
R26965 VDD.n33 VDD.n32 9.0005
R26966 VDD.n152 VDD.n151 9.0005
R26967 VDD.n30 VDD.n29 9.0005
R26968 VDD.n157 VDD.n156 9.0005
R26969 VDD.n25 VDD.n24 9.0005
R26970 VDD.n164 VDD.n163 9.0005
R26971 VDD.n22 VDD.n21 9.0005
R26972 VDD.n169 VDD.n168 9.0005
R26973 VDD.n17 VDD.n16 9.0005
R26974 VDD.n176 VDD.n175 9.0005
R26975 VDD.n14 VDD.n13 9.0005
R26976 VDD.n182 VDD.n181 9.0005
R26977 VDD.n9 VDD.n8 9.0005
R26978 VDD.n189 VDD.n188 9.0005
R26979 VDD.n190 VDD.n4 9.0005
R26980 VDD.n2015 VDD.n5 9.0005
R26981 VDD.n2014 VDD.n2013 9.0005
R26982 VDD.n6 VDD.n1 9.0005
R26983 VDD.n2040 VDD.n2039 9.0005
R26984 VDD.n80 VDD.n70 9.0005
R26985 VDD.n82 VDD.n81 9.0005
R26986 VDD.n66 VDD.n65 9.0005
R26987 VDD.n91 VDD.n90 9.0005
R26988 VDD.n92 VDD.n64 9.0005
R26989 VDD.n95 VDD.n94 9.0005
R26990 VDD.n93 VDD.n58 9.0005
R26991 VDD.n103 VDD.n57 9.0005
R26992 VDD.n105 VDD.n104 9.0005
R26993 VDD.n106 VDD.n56 9.0005
R26994 VDD.n108 VDD.n107 9.0005
R26995 VDD.n109 VDD.n55 9.0005
R26996 VDD.n111 VDD.n110 9.0005
R26997 VDD.n112 VDD.n54 9.0005
R26998 VDD.n114 VDD.n113 9.0005
R26999 VDD.n115 VDD.n53 9.0005
R27000 VDD.n117 VDD.n116 9.0005
R27001 VDD.n118 VDD.n52 9.0005
R27002 VDD.n120 VDD.n119 9.0005
R27003 VDD.n121 VDD.n51 9.0005
R27004 VDD.n123 VDD.n122 9.0005
R27005 VDD.n124 VDD.n50 9.0005
R27006 VDD.n126 VDD.n125 9.0005
R27007 VDD.n44 VDD.n43 9.0005
R27008 VDD.n135 VDD.n134 9.0005
R27009 VDD.n136 VDD.n42 9.0005
R27010 VDD.n138 VDD.n137 9.0005
R27011 VDD.n36 VDD.n35 9.0005
R27012 VDD.n147 VDD.n146 9.0005
R27013 VDD.n148 VDD.n34 9.0005
R27014 VDD.n150 VDD.n149 9.0005
R27015 VDD.n28 VDD.n27 9.0005
R27016 VDD.n159 VDD.n158 9.0005
R27017 VDD.n160 VDD.n26 9.0005
R27018 VDD.n162 VDD.n161 9.0005
R27019 VDD.n20 VDD.n19 9.0005
R27020 VDD.n171 VDD.n170 9.0005
R27021 VDD.n172 VDD.n18 9.0005
R27022 VDD.n174 VDD.n173 9.0005
R27023 VDD.n12 VDD.n11 9.0005
R27024 VDD.n184 VDD.n183 9.0005
R27025 VDD.n185 VDD.n10 9.0005
R27026 VDD.n187 VDD.n186 9.0005
R27027 VDD.n3 VDD.n2 9.0005
R27028 VDD.n2017 VDD.n2016 9.0005
R27029 VDD.n2018 VDD.n0 9.0005
R27030 VDD.n50 VDD.n49 9.0005
R27031 VDD.n127 VDD.n126 9.0005
R27032 VDD.n45 VDD.n44 9.0005
R27033 VDD.n134 VDD.n133 9.0005
R27034 VDD.n42 VDD.n41 9.0005
R27035 VDD.n139 VDD.n138 9.0005
R27036 VDD.n37 VDD.n36 9.0005
R27037 VDD.n146 VDD.n145 9.0005
R27038 VDD.n34 VDD.n33 9.0005
R27039 VDD.n151 VDD.n150 9.0005
R27040 VDD.n29 VDD.n28 9.0005
R27041 VDD.n158 VDD.n157 9.0005
R27042 VDD.n26 VDD.n25 9.0005
R27043 VDD.n163 VDD.n162 9.0005
R27044 VDD.n21 VDD.n20 9.0005
R27045 VDD.n170 VDD.n169 9.0005
R27046 VDD.n18 VDD.n17 9.0005
R27047 VDD.n175 VDD.n174 9.0005
R27048 VDD.n13 VDD.n12 9.0005
R27049 VDD.n183 VDD.n182 9.0005
R27050 VDD.n10 VDD.n9 9.0005
R27051 VDD.n188 VDD.n187 9.0005
R27052 VDD.n4 VDD.n3 9.0005
R27053 VDD.n2016 VDD.n2015 9.0005
R27054 VDD.n2014 VDD.n0 9.0005
R27055 VDD.n2054 VDD.n1 9.0005
R27056 VDD.n2054 VDD.n2053 9.0005
R27057 VDD.n84 VDD.n70 9.0005
R27058 VDD.n83 VDD.n82 9.0005
R27059 VDD.n67 VDD.n66 9.0005
R27060 VDD.n90 VDD.n89 9.0005
R27061 VDD.n64 VDD.n63 9.0005
R27062 VDD.n96 VDD.n95 9.0005
R27063 VDD.n59 VDD.n58 9.0005
R27064 VDD.n103 VDD.n102 9.0005
R27065 VDD.n83 VDD.n69 9.0005
R27066 VDD.n68 VDD.n67 9.0005
R27067 VDD.n89 VDD.n88 9.0005
R27068 VDD.n63 VDD.n62 9.0005
R27069 VDD.n97 VDD.n96 9.0005
R27070 VDD.n60 VDD.n59 9.0005
R27071 VDD.n102 VDD.n101 9.0005
R27072 VDD.n86 VDD.n68 9.0005
R27073 VDD.n88 VDD.n87 9.0005
R27074 VDD.n62 VDD.n61 9.0005
R27075 VDD.n98 VDD.n97 9.0005
R27076 VDD.n99 VDD.n60 9.0005
R27077 VDD.n101 VDD.n100 9.0005
R27078 VDD.n48 VDD.n47 9.0005
R27079 VDD.n129 VDD.n128 9.0005
R27080 VDD.n130 VDD.n46 9.0005
R27081 VDD.n132 VDD.n131 9.0005
R27082 VDD.n40 VDD.n39 9.0005
R27083 VDD.n141 VDD.n140 9.0005
R27084 VDD.n142 VDD.n38 9.0005
R27085 VDD.n144 VDD.n143 9.0005
R27086 VDD.n32 VDD.n31 9.0005
R27087 VDD.n153 VDD.n152 9.0005
R27088 VDD.n154 VDD.n30 9.0005
R27089 VDD.n156 VDD.n155 9.0005
R27090 VDD.n24 VDD.n23 9.0005
R27091 VDD.n165 VDD.n164 9.0005
R27092 VDD.n166 VDD.n22 9.0005
R27093 VDD.n168 VDD.n167 9.0005
R27094 VDD.n16 VDD.n15 9.0005
R27095 VDD.n177 VDD.n176 9.0005
R27096 VDD.n178 VDD.n14 9.0005
R27097 VDD.n181 VDD.n180 9.0005
R27098 VDD.n179 VDD.n8 9.0005
R27099 VDD.n189 VDD.n7 9.0005
R27100 VDD.n191 VDD.n190 9.0005
R27101 VDD.n192 VDD.n5 9.0005
R27102 VDD.n2013 VDD.n2012 9.0005
R27103 VDD.n2011 VDD.n6 9.0005
R27104 VDD.n2010 VDD.n2009 9.0005
R27105 VDD.n2008 VDD.n193 9.0005
R27106 VDD.n2007 VDD.n2006 9.0005
R27107 VDD.n2005 VDD.n197 9.0005
R27108 VDD.n2004 VDD.n2003 9.0005
R27109 VDD.n2002 VDD.n198 9.0005
R27110 VDD.n2001 VDD.n2000 9.0005
R27111 VDD.n1999 VDD.n202 9.0005
R27112 VDD.n1998 VDD.n1997 9.0005
R27113 VDD.n1996 VDD.n203 9.0005
R27114 VDD.n1995 VDD.n1994 9.0005
R27115 VDD.n1993 VDD.n207 9.0005
R27116 VDD.n1992 VDD.n1991 9.0005
R27117 VDD.n1990 VDD.n208 9.0005
R27118 VDD.n1989 VDD.n1988 9.0005
R27119 VDD.n1987 VDD.n212 9.0005
R27120 VDD.n1986 VDD.n1985 9.0005
R27121 VDD.n1984 VDD.n213 9.0005
R27122 VDD.n1983 VDD.n1982 9.0005
R27123 VDD.n1981 VDD.n217 9.0005
R27124 VDD.n1980 VDD.n1979 9.0005
R27125 VDD.n1978 VDD.n218 9.0005
R27126 VDD.n1977 VDD.n1976 9.0005
R27127 VDD.n1975 VDD.n222 9.0005
R27128 VDD.n1974 VDD.n1973 9.0005
R27129 VDD.n1972 VDD.n223 9.0005
R27130 VDD.n1971 VDD.n1970 9.0005
R27131 VDD.n1969 VDD.n227 9.0005
R27132 VDD.n1968 VDD.n1967 9.0005
R27133 VDD.n1966 VDD.n228 9.0005
R27134 VDD.n1965 VDD.n1964 9.0005
R27135 VDD.n1963 VDD.n232 9.0005
R27136 VDD.n1962 VDD.n1961 9.0005
R27137 VDD.n1960 VDD.n233 9.0005
R27138 VDD.n1959 VDD.n1958 9.0005
R27139 VDD.n1957 VDD.n237 9.0005
R27140 VDD.n1956 VDD.n1955 9.0005
R27141 VDD.n1954 VDD.n238 9.0005
R27142 VDD.n1953 VDD.n1952 9.0005
R27143 VDD.n1951 VDD.n242 9.0005
R27144 VDD.n1950 VDD.n1949 9.0005
R27145 VDD.n1948 VDD.n243 9.0005
R27146 VDD.n1947 VDD.n1946 9.0005
R27147 VDD.n1945 VDD.n247 9.0005
R27148 VDD.n1944 VDD.n1943 9.0005
R27149 VDD.n1942 VDD.n248 9.0005
R27150 VDD.n1941 VDD.n1940 9.0005
R27151 VDD.n2046 VDD.n2045 8.5005
R27152 VDD.n2036 VDD.n2034 8.5005
R27153 VDD.n2050 VDD.n2019 8.5005
R27154 VDD.n72 VDD.n71 8.47111
R27155 VDD.n307 VDD.n287 7.96796
R27156 VDD.n308 VDD.n307 7.9321
R27157 VDD.n2048 VDD.n2021 7.9321
R27158 VDD.n2049 VDD.n2048 7.9321
R27159 VDD.n1940 VDD.n1939 6.82903
R27160 VDD.n307 VDD.n306 6.0367
R27161 VDD.n2048 VDD.n2047 6.0005
R27162 VDD.n299 VDD.n296 5.65698
R27163 VDD.n310 VDD.n285 5.65698
R27164 VDD.n2045 VDD.n2044 5.65698
R27165 VDD.n2036 VDD.n2035 5.65698
R27166 VDD.n2025 VDD.n2019 5.65698
R27167 VDD.n305 VDD.n291 5.65698
R27168 VDD.n254 VDD.n252 5.61485
R27169 VDD.n311 VDD.n310 5.61485
R27170 VDD.n77 VDD.n71 5.61485
R27171 VDD.n310 VDD.n309 5.61447
R27172 VDD.n556 VDD.n551 4.70565
R27173 VDD.n570 VDD.n569 4.6277
R27174 VDD.n576 VDD.n566 4.597
R27175 VDD.n86 VDD.n85 4.56021
R27176 VDD.n582 VDD.n581 4.5005
R27177 VDD.n522 VDD.n521 4.46912
R27178 VDD.n443 VDD.n442 4.4685
R27179 VDD.n310 VDD.n286 4.24021
R27180 VDD.n2052 VDD.n2019 4.18639
R27181 VDD.n256 VDD.n252 4.17719
R27182 VDD.n79 VDD.n71 4.17719
R27183 VDD.n76 VDD.n71 4.17719
R27184 VDD.n2045 VDD.n2022 3.38382
R27185 VDD.n2036 VDD.n2033 3.38382
R27186 VDD.n2020 VDD.n2019 3.38382
R27187 VDD.n2011 VDD.n2010 2.93984
R27188 VDD.n299 VDD.n287 2.81935
R27189 VDD.n306 VDD.n305 2.81935
R27190 VDD.n305 VDD.n288 2.35437
R27191 VDD.n300 VDD.n299 2.35437
R27192 VDD.n310 VDD.n281 2.35437
R27193 VDD.n2024 VDD.n2019 2.35393
R27194 VDD.n2036 VDD.n2030 2.35371
R27195 VDD.n253 VDD.n252 2.29824
R27196 VDD.n1463 VDD.n1462 2.2505
R27197 VDD.n1442 VDD.n1441 2.2505
R27198 VDD.n1437 VDD.n918 2.2505
R27199 VDD.n1435 VDD.n920 2.2505
R27200 VDD.n1431 VDD.n923 2.2505
R27201 VDD.n1429 VDD.n925 2.2505
R27202 VDD.n1425 VDD.n928 2.2505
R27203 VDD.n1423 VDD.n930 2.2505
R27204 VDD.n994 VDD.n931 2.2505
R27205 VDD.n1418 VDD.n934 2.2505
R27206 VDD.n1197 VDD.n936 2.2505
R27207 VDD.n1412 VDD.n939 2.2505
R27208 VDD.n1244 VDD.n941 2.2505
R27209 VDD.n1406 VDD.n944 2.2505
R27210 VDD.n1276 VDD.n946 2.2505
R27211 VDD.n1851 VDD.n1847 2.2505
R27212 VDD.n1845 VDD.n1844 2.2505
R27213 VDD.n1824 VDD.n1823 2.2505
R27214 VDD.n1821 VDD.n1820 2.2505
R27215 VDD.n1795 VDD.n1794 2.2505
R27216 VDD.n1792 VDD.n1791 2.2505
R27217 VDD.n1775 VDD.n1774 2.2505
R27218 VDD.n1773 VDD.n712 2.2505
R27219 VDD.n714 VDD.n713 2.2505
R27220 VDD.n1745 VDD.n723 2.2505
R27221 VDD.n725 VDD.n724 2.2505
R27222 VDD.n1720 VDD.n736 2.2505
R27223 VDD.n738 VDD.n737 2.2505
R27224 VDD.n1700 VDD.n748 2.2505
R27225 VDD.n750 VDD.n749 2.2505
R27226 VDD.n1852 VDD.n1851 2.2505
R27227 VDD.n1844 VDD.n1843 2.2505
R27228 VDD.n1825 VDD.n1824 2.2505
R27229 VDD.n1820 VDD.n1819 2.2505
R27230 VDD.n1796 VDD.n1795 2.2505
R27231 VDD.n1791 VDD.n1790 2.2505
R27232 VDD.n1776 VDD.n1775 2.2505
R27233 VDD.n1764 VDD.n712 2.2505
R27234 VDD.n1755 VDD.n714 2.2505
R27235 VDD.n727 VDD.n723 2.2505
R27236 VDD.n1731 VDD.n725 2.2505
R27237 VDD.n740 VDD.n736 2.2505
R27238 VDD.n1706 VDD.n738 2.2505
R27239 VDD.n758 VDD.n748 2.2505
R27240 VDD.n1687 VDD.n750 2.2505
R27241 VDD.n1469 VDD.n1468 2.2505
R27242 VDD.n878 VDD.n870 2.2505
R27243 VDD.n1481 VDD.n866 2.2505
R27244 VDD.n1490 VDD.n1489 2.2505
R27245 VDD.n868 VDD.n864 2.2505
R27246 VDD.n1495 VDD.n1494 2.2505
R27247 VDD.n1505 VDD.n852 2.2505
R27248 VDD.n1514 VDD.n1513 2.2505
R27249 VDD.n849 VDD.n845 2.2505
R27250 VDD.n1526 VDD.n1525 2.2505
R27251 VDD.n850 VDD.n838 2.2505
R27252 VDD.n1521 VDD.n836 2.2505
R27253 VDD.n1520 VDD.n834 2.2505
R27254 VDD.n1519 VDD.n832 2.2505
R27255 VDD.n1552 VDD.n823 2.2505
R27256 VDD.n1570 VDD.n1569 2.2505
R27257 VDD.n1562 VDD.n821 2.2505
R27258 VDD.n1575 VDD.n1574 2.2505
R27259 VDD.n1578 VDD.n810 2.2505
R27260 VDD.n1594 VDD.n1593 2.2505
R27261 VDD.n812 VDD.n808 2.2505
R27262 VDD.n1599 VDD.n1598 2.2505
R27263 VDD.n1603 VDD.n797 2.2505
R27264 VDD.n1620 VDD.n1619 2.2505
R27265 VDD.n1611 VDD.n795 2.2505
R27266 VDD.n1625 VDD.n1624 2.2505
R27267 VDD.n1628 VDD.n784 2.2505
R27268 VDD.n1646 VDD.n1645 2.2505
R27269 VDD.n1638 VDD.n781 2.2505
R27270 VDD.n1652 VDD.n1651 2.2505
R27271 VDD.n782 VDD.n776 2.2505
R27272 VDD.n1666 VDD.n768 2.2505
R27273 VDD.n1680 VDD.n1679 2.2505
R27274 VDD.n766 VDD.n763 2.2505
R27275 VDD.n1682 VDD.n766 2.2505
R27276 VDD.n1681 VDD.n1680 2.2505
R27277 VDD.n768 VDD.n767 2.2505
R27278 VDD.n1649 VDD.n782 2.2505
R27279 VDD.n1651 VDD.n1650 2.2505
R27280 VDD.n1648 VDD.n781 2.2505
R27281 VDD.n1647 VDD.n1646 2.2505
R27282 VDD.n784 VDD.n783 2.2505
R27283 VDD.n1624 VDD.n1623 2.2505
R27284 VDD.n1622 VDD.n795 2.2505
R27285 VDD.n1621 VDD.n1620 2.2505
R27286 VDD.n797 VDD.n796 2.2505
R27287 VDD.n1598 VDD.n1597 2.2505
R27288 VDD.n1596 VDD.n808 2.2505
R27289 VDD.n1595 VDD.n1594 2.2505
R27290 VDD.n810 VDD.n809 2.2505
R27291 VDD.n1574 VDD.n1573 2.2505
R27292 VDD.n1572 VDD.n821 2.2505
R27293 VDD.n1571 VDD.n1570 2.2505
R27294 VDD.n823 VDD.n822 2.2505
R27295 VDD.n1519 VDD.n1518 2.2505
R27296 VDD.n1520 VDD.n1517 2.2505
R27297 VDD.n1522 VDD.n1521 2.2505
R27298 VDD.n1523 VDD.n850 2.2505
R27299 VDD.n1525 VDD.n1524 2.2505
R27300 VDD.n1516 VDD.n849 2.2505
R27301 VDD.n1515 VDD.n1514 2.2505
R27302 VDD.n852 VDD.n851 2.2505
R27303 VDD.n1494 VDD.n1493 2.2505
R27304 VDD.n1492 VDD.n864 2.2505
R27305 VDD.n1491 VDD.n1490 2.2505
R27306 VDD.n866 VDD.n865 2.2505
R27307 VDD.n1466 VDD.n878 2.2505
R27308 VDD.n1468 VDD.n1467 2.2505
R27309 VDD.n1464 VDD.n1463 2.2505
R27310 VDD.n1441 VDD.n1440 2.2505
R27311 VDD.n1438 VDD.n1437 2.2505
R27312 VDD.n1435 VDD.n1434 2.2505
R27313 VDD.n1432 VDD.n1431 2.2505
R27314 VDD.n1429 VDD.n1428 2.2505
R27315 VDD.n1426 VDD.n1425 2.2505
R27316 VDD.n1423 VDD.n1422 2.2505
R27317 VDD.n1421 VDD.n931 2.2505
R27318 VDD.n1418 VDD.n932 2.2505
R27319 VDD.n1415 VDD.n936 2.2505
R27320 VDD.n1412 VDD.n937 2.2505
R27321 VDD.n1409 VDD.n941 2.2505
R27322 VDD.n1406 VDD.n942 2.2505
R27323 VDD.n1403 VDD.n946 2.2505
R27324 VDD.n1848 VDD.n667 2.2505
R27325 VDD.n1875 VDD.n666 2.2505
R27326 VDD.n1876 VDD.n665 2.2505
R27327 VDD.n664 VDD.n658 2.2505
R27328 VDD.n663 VDD.n662 2.2505
R27329 VDD.n661 VDD.n660 2.2505
R27330 VDD.n659 VDD.n642 2.2505
R27331 VDD.n1897 VDD.n641 2.2505
R27332 VDD.n1898 VDD.n640 2.2505
R27333 VDD.n639 VDD.n637 2.2505
R27334 VDD.n638 VDD.n622 2.2505
R27335 VDD.n1910 VDD.n621 2.2505
R27336 VDD.n1911 VDD.n620 2.2505
R27337 VDD.n619 VDD.n617 2.2505
R27338 VDD.n618 VDD.n602 2.2505
R27339 VDD.n1922 VDD.n601 2.2505
R27340 VDD.n1923 VDD.n600 2.2505
R27341 VDD.n1345 VDD.n599 2.2505
R27342 VDD.n1347 VDD.n1346 2.2505
R27343 VDD.n1349 VDD.n1348 2.2505
R27344 VDD.n1351 VDD.n1350 2.2505
R27345 VDD.n1353 VDD.n1352 2.2505
R27346 VDD.n1355 VDD.n1354 2.2505
R27347 VDD.n1357 VDD.n1356 2.2505
R27348 VDD.n1358 VDD.n1344 2.2505
R27349 VDD.n1343 VDD.n1328 2.2505
R27350 VDD.n1370 VDD.n1327 2.2505
R27351 VDD.n1371 VDD.n1326 2.2505
R27352 VDD.n1325 VDD.n1312 2.2505
R27353 VDD.n1382 VDD.n1311 2.2505
R27354 VDD.n1383 VDD.n1310 2.2505
R27355 VDD.n1309 VDD.n1306 2.2505
R27356 VDD.n1308 VDD.n1307 2.2505
R27357 VDD.n948 VDD.n947 2.2505
R27358 VDD.n1298 VDD.n948 2.2505
R27359 VDD.n1307 VDD.n1302 2.2505
R27360 VDD.n1306 VDD.n1303 2.2505
R27361 VDD.n1384 VDD.n1383 2.2505
R27362 VDD.n1382 VDD.n1381 2.2505
R27363 VDD.n1322 VDD.n1312 2.2505
R27364 VDD.n1372 VDD.n1371 2.2505
R27365 VDD.n1370 VDD.n1369 2.2505
R27366 VDD.n1340 VDD.n1328 2.2505
R27367 VDD.n1359 VDD.n1358 2.2505
R27368 VDD.n599 VDD.n584 2.2505
R27369 VDD.n1924 VDD.n1923 2.2505
R27370 VDD.n1922 VDD.n1921 2.2505
R27371 VDD.n611 VDD.n602 2.2505
R27372 VDD.n617 VDD.n615 2.2505
R27373 VDD.n1912 VDD.n1911 2.2505
R27374 VDD.n1910 VDD.n1909 2.2505
R27375 VDD.n631 VDD.n622 2.2505
R27376 VDD.n637 VDD.n635 2.2505
R27377 VDD.n1899 VDD.n1898 2.2505
R27378 VDD.n1897 VDD.n1896 2.2505
R27379 VDD.n650 VDD.n642 2.2505
R27380 VDD.n661 VDD.n651 2.2505
R27381 VDD.n662 VDD.n653 2.2505
R27382 VDD.n658 VDD.n655 2.2505
R27383 VDD.n1877 VDD.n1876 2.2505
R27384 VDD.n1875 VDD.n1874 2.2505
R27385 VDD.n672 VDD.n667 2.2505
R27386 VDD.n1286 VDD.n949 2.2005
R27387 VDD.n1277 VDD.n956 2.2005
R27388 VDD.n1279 VDD.n1278 2.2005
R27389 VDD.n1270 VDD.n1269 2.2005
R27390 VDD.n1268 VDD.n1267 2.2005
R27391 VDD.n1262 VDD.n961 2.2005
R27392 VDD.n1253 VDD.n964 2.2005
R27393 VDD.n1255 VDD.n1254 2.2005
R27394 VDD.n1245 VDD.n966 2.2005
R27395 VDD.n1247 VDD.n1246 2.2005
R27396 VDD.n1243 VDD.n1242 2.2005
R27397 VDD.n1235 VDD.n969 2.2005
R27398 VDD.n1229 VDD.n1228 2.2005
R27399 VDD.n1227 VDD.n1226 2.2005
R27400 VDD.n1222 VDD.n1221 2.2005
R27401 VDD.n1220 VDD.n1219 2.2005
R27402 VDD.n1214 VDD.n1213 2.2005
R27403 VDD.n1212 VDD.n1211 2.2005
R27404 VDD.n1205 VDD.n981 2.2005
R27405 VDD.n1199 VDD.n1198 2.2005
R27406 VDD.n1196 VDD.n1195 2.2005
R27407 VDD.n1186 VDD.n986 2.2005
R27408 VDD.n1188 VDD.n1187 2.2005
R27409 VDD.n1181 VDD.n1180 2.2005
R27410 VDD.n1179 VDD.n1178 2.2005
R27411 VDD.n1172 VDD.n1171 2.2005
R27412 VDD.n1170 VDD.n1169 2.2005
R27413 VDD.n1163 VDD.n1162 2.2005
R27414 VDD.n1161 VDD.n1160 2.2005
R27415 VDD.n1154 VDD.n1153 2.2005
R27416 VDD.n1152 VDD.n1151 2.2005
R27417 VDD.n1145 VDD.n1144 2.2005
R27418 VDD.n1143 VDD.n1142 2.2005
R27419 VDD.n1137 VDD.n1005 2.2005
R27420 VDD.n1128 VDD.n1009 2.2005
R27421 VDD.n1130 VDD.n1129 2.2005
R27422 VDD.n1126 VDD.n1125 2.2005
R27423 VDD.n1118 VDD.n1012 2.2005
R27424 VDD.n1112 VDD.n1111 2.2005
R27425 VDD.n1110 VDD.n1109 2.2005
R27426 VDD.n1105 VDD.n1104 2.2005
R27427 VDD.n1103 VDD.n1102 2.2005
R27428 VDD.n1097 VDD.n1096 2.2005
R27429 VDD.n1095 VDD.n1094 2.2005
R27430 VDD.n1088 VDD.n1024 2.2005
R27431 VDD.n1082 VDD.n1081 2.2005
R27432 VDD.n1079 VDD.n1078 2.2005
R27433 VDD.n1069 VDD.n1029 2.2005
R27434 VDD.n1071 VDD.n1070 2.2005
R27435 VDD.n1064 VDD.n1063 2.2005
R27436 VDD.n1062 VDD.n1061 2.2005
R27437 VDD.n1055 VDD.n1054 2.2005
R27438 VDD.n1053 VDD.n1052 2.2005
R27439 VDD.n1046 VDD.n1045 2.2005
R27440 VDD.n1043 VDD.n915 2.2005
R27441 VDD.n1444 VDD.n1443 2.2005
R27442 VDD.n1449 VDD.n911 2.2005
R27443 VDD.n910 VDD.n907 2.2005
R27444 VDD.n1456 VDD.n882 2.2005
R27445 VDD.n1461 VDD.n1460 2.2005
R27446 VDD.n902 VDD.n881 2.2005
R27447 VDD.n679 VDD.n671 2.2005
R27448 VDD.n1686 VDD.n762 2.2005
R27449 VDD.n1689 VDD.n1688 2.2005
R27450 VDD.n753 VDD.n751 2.2005
R27451 VDD.n1696 VDD.n1695 2.2005
R27452 VDD.n1694 VDD.n752 2.2005
R27453 VDD.n760 VDD.n759 2.2005
R27454 VDD.n757 VDD.n756 2.2005
R27455 VDD.n754 VDD.n747 2.2005
R27456 VDD.n1704 VDD.n744 2.2005
R27457 VDD.n1708 VDD.n1707 2.2005
R27458 VDD.n1705 VDD.n746 2.2005
R27459 VDD.n745 VDD.n739 2.2005
R27460 VDD.n1716 VDD.n1715 2.2005
R27461 VDD.n1714 VDD.n741 2.2005
R27462 VDD.n735 VDD.n734 2.2005
R27463 VDD.n1725 VDD.n1724 2.2005
R27464 VDD.n1727 VDD.n733 2.2005
R27465 VDD.n1729 VDD.n1728 2.2005
R27466 VDD.n1730 VDD.n731 2.2005
R27467 VDD.n1733 VDD.n1732 2.2005
R27468 VDD.n732 VDD.n726 2.2005
R27469 VDD.n1741 VDD.n1740 2.2005
R27470 VDD.n1739 VDD.n728 2.2005
R27471 VDD.n722 VDD.n721 2.2005
R27472 VDD.n1750 VDD.n1749 2.2005
R27473 VDD.n1751 VDD.n720 2.2005
R27474 VDD.n1754 VDD.n1753 2.2005
R27475 VDD.n1756 VDD.n719 2.2005
R27476 VDD.n1758 VDD.n1757 2.2005
R27477 VDD.n717 VDD.n715 2.2005
R27478 VDD.n1769 VDD.n1768 2.2005
R27479 VDD.n1767 VDD.n716 2.2005
R27480 VDD.n1766 VDD.n1765 2.2005
R27481 VDD.n1762 VDD.n711 2.2005
R27482 VDD.n1777 VDD.n708 2.2005
R27483 VDD.n1781 VDD.n1780 2.2005
R27484 VDD.n1778 VDD.n710 2.2005
R27485 VDD.n709 VDD.n703 2.2005
R27486 VDD.n1789 VDD.n1788 2.2005
R27487 VDD.n1787 VDD.n705 2.2005
R27488 VDD.n699 VDD.n698 2.2005
R27489 VDD.n1798 VDD.n1797 2.2005
R27490 VDD.n1800 VDD.n697 2.2005
R27491 VDD.n1802 VDD.n1801 2.2005
R27492 VDD.n1803 VDD.n696 2.2005
R27493 VDD.n1806 VDD.n1805 2.2005
R27494 VDD.n694 VDD.n692 2.2005
R27495 VDD.n1818 VDD.n1817 2.2005
R27496 VDD.n1816 VDD.n693 2.2005
R27497 VDD.n1814 VDD.n1813 2.2005
R27498 VDD.n1811 VDD.n688 2.2005
R27499 VDD.n1826 VDD.n687 2.2005
R27500 VDD.n1830 VDD.n1829 2.2005
R27501 VDD.n1827 VDD.n685 2.2005
R27502 VDD.n1835 VDD.n683 2.2005
R27503 VDD.n1842 VDD.n1841 2.2005
R27504 VDD.n1839 VDD.n684 2.2005
R27505 VDD.n1838 VDD.n1837 2.2005
R27506 VDD.n678 VDD.n677 2.2005
R27507 VDD.n1854 VDD.n1853 2.2005
R27508 VDD.n1294 VDD.n950 2.2005
R27509 VDD.n1299 VDD.n1296 2.2005
R27510 VDD.n1392 VDD.n1300 2.2005
R27511 VDD.n1391 VDD.n1390 2.2005
R27512 VDD.n1389 VDD.n1388 2.2005
R27513 VDD.n1387 VDD.n1386 2.2005
R27514 VDD.n1385 VDD.n1304 2.2005
R27515 VDD.n1314 VDD.n1305 2.2005
R27516 VDD.n1380 VDD.n1379 2.2005
R27517 VDD.n1315 VDD.n1313 2.2005
R27518 VDD.n1323 VDD.n1320 2.2005
R27519 VDD.n1374 VDD.n1373 2.2005
R27520 VDD.n1324 VDD.n1321 2.2005
R27521 VDD.n1331 VDD.n1329 2.2005
R27522 VDD.n1368 VDD.n1367 2.2005
R27523 VDD.n1366 VDD.n1330 2.2005
R27524 VDD.n1341 VDD.n1333 2.2005
R27525 VDD.n1342 VDD.n1338 2.2005
R27526 VDD.n1361 VDD.n1360 2.2005
R27527 VDD.n1339 VDD.n583 2.2005
R27528 VDD.n1927 VDD.n596 2.2005
R27529 VDD.n1926 VDD.n1925 2.2005
R27530 VDD.n598 VDD.n597 2.2005
R27531 VDD.n606 VDD.n603 2.2005
R27532 VDD.n1920 VDD.n1919 2.2005
R27533 VDD.n607 VDD.n604 2.2005
R27534 VDD.n613 VDD.n612 2.2005
R27535 VDD.n614 VDD.n609 2.2005
R27536 VDD.n1914 VDD.n1913 2.2005
R27537 VDD.n616 VDD.n610 2.2005
R27538 VDD.n626 VDD.n623 2.2005
R27539 VDD.n1908 VDD.n1907 2.2005
R27540 VDD.n627 VDD.n624 2.2005
R27541 VDD.n633 VDD.n632 2.2005
R27542 VDD.n634 VDD.n629 2.2005
R27543 VDD.n1902 VDD.n1901 2.2005
R27544 VDD.n1900 VDD.n630 2.2005
R27545 VDD.n646 VDD.n636 2.2005
R27546 VDD.n647 VDD.n643 2.2005
R27547 VDD.n1895 VDD.n1894 2.2005
R27548 VDD.n1893 VDD.n644 2.2005
R27549 VDD.n1892 VDD.n1891 2.2005
R27550 VDD.n1890 VDD.n1889 2.2005
R27551 VDD.n1888 VDD.n1887 2.2005
R27552 VDD.n1886 VDD.n1885 2.2005
R27553 VDD.n1884 VDD.n1883 2.2005
R27554 VDD.n1882 VDD.n1881 2.2005
R27555 VDD.n1880 VDD.n1879 2.2005
R27556 VDD.n1878 VDD.n656 2.2005
R27557 VDD.n1865 VDD.n657 2.2005
R27558 VDD.n1864 VDD.n668 2.2005
R27559 VDD.n1873 VDD.n1872 2.2005
R27560 VDD.n1871 VDD.n669 2.2005
R27561 VDD.n890 VDD.n876 2.2005
R27562 VDD.n1470 VDD.n875 2.2005
R27563 VDD.n1472 VDD.n1471 2.2005
R27564 VDD.n1479 VDD.n1478 2.2005
R27565 VDD.n1480 VDD.n869 2.2005
R27566 VDD.n1483 VDD.n1482 2.2005
R27567 VDD.n1485 VDD.n867 2.2005
R27568 VDD.n1488 VDD.n1487 2.2005
R27569 VDD.n863 VDD.n861 2.2005
R27570 VDD.n1497 VDD.n1496 2.2005
R27571 VDD.n857 VDD.n856 2.2005
R27572 VDD.n1504 VDD.n1503 2.2005
R27573 VDD.n1507 VDD.n1506 2.2005
R27574 VDD.n1509 VDD.n853 2.2005
R27575 VDD.n1512 VDD.n1511 2.2005
R27576 VDD.n854 VDD.n843 2.2005
R27577 VDD.n1529 VDD.n1528 2.2005
R27578 VDD.n1527 VDD.n844 2.2005
R27579 VDD.n848 VDD.n847 2.2005
R27580 VDD.n846 VDD.n839 2.2005
R27581 VDD.n1537 VDD.n1536 2.2005
R27582 VDD.n1539 VDD.n1538 2.2005
R27583 VDD.n1541 VDD.n1540 2.2005
R27584 VDD.n1543 VDD.n1542 2.2005
R27585 VDD.n1545 VDD.n1544 2.2005
R27586 VDD.n1547 VDD.n1546 2.2005
R27587 VDD.n1550 VDD.n1549 2.2005
R27588 VDD.n1551 VDD.n830 2.2005
R27589 VDD.n1554 VDD.n1553 2.2005
R27590 VDD.n826 VDD.n824 2.2005
R27591 VDD.n1568 VDD.n1567 2.2005
R27592 VDD.n1566 VDD.n825 2.2005
R27593 VDD.n1564 VDD.n1563 2.2005
R27594 VDD.n1560 VDD.n820 2.2005
R27595 VDD.n1576 VDD.n818 2.2005
R27596 VDD.n1580 VDD.n1579 2.2005
R27597 VDD.n1577 VDD.n814 2.2005
R27598 VDD.n1586 VDD.n811 2.2005
R27599 VDD.n1592 VDD.n1591 2.2005
R27600 VDD.n1589 VDD.n813 2.2005
R27601 VDD.n1587 VDD.n807 2.2005
R27602 VDD.n1600 VDD.n805 2.2005
R27603 VDD.n1605 VDD.n1604 2.2005
R27604 VDD.n1602 VDD.n1601 2.2005
R27605 VDD.n800 VDD.n798 2.2005
R27606 VDD.n1618 VDD.n1617 2.2005
R27607 VDD.n1615 VDD.n799 2.2005
R27608 VDD.n1613 VDD.n1612 2.2005
R27609 VDD.n794 VDD.n792 2.2005
R27610 VDD.n1631 VDD.n1630 2.2005
R27611 VDD.n1629 VDD.n793 2.2005
R27612 VDD.n1627 VDD.n1626 2.2005
R27613 VDD.n789 VDD.n785 2.2005
R27614 VDD.n1644 VDD.n1643 2.2005
R27615 VDD.n1641 VDD.n786 2.2005
R27616 VDD.n1640 VDD.n1639 2.2005
R27617 VDD.n780 VDD.n779 2.2005
R27618 VDD.n1655 VDD.n1654 2.2005
R27619 VDD.n1653 VDD.n777 2.2005
R27620 VDD.n1664 VDD.n1663 2.2005
R27621 VDD.n1668 VDD.n1667 2.2005
R27622 VDD.n1665 VDD.n773 2.2005
R27623 VDD.n772 VDD.n769 2.2005
R27624 VDD.n1678 VDD.n1677 2.2005
R27625 VDD.n1676 VDD.n770 2.2005
R27626 VDD.n1934 VDD.n587 2.2005
R27627 VDD.n909 VDD.n880 1.8005
R27628 VDD.n1037 VDD.n916 1.8005
R27629 VDD.n1436 VDD.n919 1.8005
R27630 VDD.n1080 VDD.n921 1.8005
R27631 VDD.n1430 VDD.n924 1.8005
R27632 VDD.n1127 VDD.n926 1.8005
R27633 VDD.n1424 VDD.n929 1.8005
R27634 VDD.n1419 VDD.n933 1.8005
R27635 VDD.n1417 VDD.n935 1.8005
R27636 VDD.n1413 VDD.n938 1.8005
R27637 VDD.n1411 VDD.n940 1.8005
R27638 VDD.n1407 VDD.n943 1.8005
R27639 VDD.n1405 VDD.n945 1.8005
R27640 VDD.n1846 VDD.n680 1.8005
R27641 VDD.n682 VDD.n681 1.8005
R27642 VDD.n1822 VDD.n689 1.8005
R27643 VDD.n691 VDD.n690 1.8005
R27644 VDD.n1793 VDD.n700 1.8005
R27645 VDD.n702 VDD.n701 1.8005
R27646 VDD.n1772 VDD.n1771 1.8005
R27647 VDD.n1747 VDD.n1746 1.8005
R27648 VDD.n1744 VDD.n1743 1.8005
R27649 VDD.n1722 VDD.n1721 1.8005
R27650 VDD.n1719 VDD.n1718 1.8005
R27651 VDD.n1702 VDD.n1701 1.8005
R27652 VDD.n1699 VDD.n1698 1.8005
R27653 VDD.n1836 VDD.n680 1.8005
R27654 VDD.n1828 VDD.n682 1.8005
R27655 VDD.n1812 VDD.n689 1.8005
R27656 VDD.n1804 VDD.n691 1.8005
R27657 VDD.n704 VDD.n700 1.8005
R27658 VDD.n1779 VDD.n702 1.8005
R27659 VDD.n1771 VDD.n1770 1.8005
R27660 VDD.n1748 VDD.n1747 1.8005
R27661 VDD.n1743 VDD.n1742 1.8005
R27662 VDD.n1723 VDD.n1722 1.8005
R27663 VDD.n1718 VDD.n1717 1.8005
R27664 VDD.n1703 VDD.n1702 1.8005
R27665 VDD.n1698 VDD.n1697 1.8005
R27666 VDD.n1685 VDD.n1684 1.8005
R27667 VDD.n1684 VDD.n1683 1.8005
R27668 VDD.n880 VDD.n879 1.8005
R27669 VDD.n1439 VDD.n916 1.8005
R27670 VDD.n1436 VDD.n917 1.8005
R27671 VDD.n1433 VDD.n921 1.8005
R27672 VDD.n1430 VDD.n922 1.8005
R27673 VDD.n1427 VDD.n926 1.8005
R27674 VDD.n1424 VDD.n927 1.8005
R27675 VDD.n1420 VDD.n1419 1.8005
R27676 VDD.n1417 VDD.n1416 1.8005
R27677 VDD.n1414 VDD.n1413 1.8005
R27678 VDD.n1411 VDD.n1410 1.8005
R27679 VDD.n1408 VDD.n1407 1.8005
R27680 VDD.n1405 VDD.n1404 1.8005
R27681 VDD.n1850 VDD.n1849 1.8005
R27682 VDD.n1850 VDD.n673 1.8005
R27683 VDD.n1935 VDD.n582 1.68488
R27684 VDD.n313 VDD.n311 1.68224
R27685 VDD.n2053 VDD 1.50225
R27686 VDD.n886 VDD.n877 1.5005
R27687 VDD.n1465 VDD.n877 1.5005
R27688 VDD.n1402 VDD.n1401 1.5005
R27689 VDD.n1401 VDD.n1400 1.5005
R27690 VDD VDD.n255 1.29335
R27691 VDD VDD.n78 1.29335
R27692 VDD VDD.n2019 1.18432
R27693 VDD.n2036 VDD 1.18273
R27694 VDD.n255 VDD 1.14327
R27695 VDD.n78 VDD 1.14327
R27696 VDD.n1934 VDD.n590 1.11718
R27697 VDD.n1934 VDD.n589 1.11718
R27698 VDD.n1934 VDD.n588 1.11718
R27699 VDD.n1396 VDD.n1295 1.1125
R27700 VDD.n1660 VDD.n775 1.10836
R27701 VDD.n1662 VDD.n1661 1.10443
R27702 VDD.n1675 VDD.n1674 1.10381
R27703 VDD.n1397 VDD.n953 1.10372
R27704 VDD.n1656 VDD.n778 1.10339
R27705 VDD.n1671 VDD.n773 1.10272
R27706 VDD.n1668 VDD.n774 1.10272
R27707 VDD.n1659 VDD.n777 1.10272
R27708 VDD.n1395 VDD.n1296 1.10263
R27709 VDD.n1392 VDD.n1297 1.10263
R27710 VDD.n1856 VDD.n1855 1.1005
R27711 VDD.n1691 VDD.n1690 1.1005
R27712 VDD.n1693 VDD.n1692 1.1005
R27713 VDD.n755 VDD.n743 1.1005
R27714 VDD.n1710 VDD.n1709 1.1005
R27715 VDD.n1711 VDD.n742 1.1005
R27716 VDD.n1713 VDD.n1712 1.1005
R27717 VDD.n1726 VDD.n730 1.1005
R27718 VDD.n1735 VDD.n1734 1.1005
R27719 VDD.n1736 VDD.n729 1.1005
R27720 VDD.n1738 VDD.n1737 1.1005
R27721 VDD.n1752 VDD.n718 1.1005
R27722 VDD.n1760 VDD.n1759 1.1005
R27723 VDD.n1768 VDD.n1761 1.1005
R27724 VDD.n1763 VDD.n707 1.1005
R27725 VDD.n1783 VDD.n1782 1.1005
R27726 VDD.n1784 VDD.n706 1.1005
R27727 VDD.n1786 VDD.n1785 1.1005
R27728 VDD.n1799 VDD.n695 1.1005
R27729 VDD.n1808 VDD.n1807 1.1005
R27730 VDD.n1810 VDD.n1809 1.1005
R27731 VDD.n1815 VDD.n686 1.1005
R27732 VDD.n1832 VDD.n1831 1.1005
R27733 VDD.n1834 VDD.n1833 1.1005
R27734 VDD.n1840 VDD.n676 1.1005
R27735 VDD.n764 VDD.n761 1.1005
R27736 VDD.n675 VDD.n674 1.1005
R27737 VDD.n1859 VDD.n1858 1.1005
R27738 VDD.n1858 VDD.n1857 1.1005
R27739 VDD.n1870 VDD.n1869 1.1005
R27740 VDD.n1868 VDD.n670 1.1005
R27741 VDD.n1867 VDD.n1866 1.1005
R27742 VDD.n1863 VDD.n654 1.1005
R27743 VDD.n1862 VDD.n652 1.1005
R27744 VDD.n1861 VDD.n649 1.1005
R27745 VDD.n1860 VDD.n648 1.1005
R27746 VDD.n645 VDD.n628 1.1005
R27747 VDD.n1904 VDD.n1903 1.1005
R27748 VDD.n1906 VDD.n1905 1.1005
R27749 VDD.n625 VDD.n608 1.1005
R27750 VDD.n1916 VDD.n1915 1.1005
R27751 VDD.n1918 VDD.n1917 1.1005
R27752 VDD.n605 VDD.n595 1.1005
R27753 VDD.n1928 VDD.n1927 1.1005
R27754 VDD.n1930 VDD.n1929 1.1005
R27755 VDD.n1932 VDD.n1931 1.1005
R27756 VDD.n594 VDD.n593 1.1005
R27757 VDD.n1335 VDD.n1334 1.1005
R27758 VDD.n1337 VDD.n1336 1.1005
R27759 VDD.n1363 VDD.n1362 1.1005
R27760 VDD.n1365 VDD.n1364 1.1005
R27761 VDD.n1332 VDD.n1319 1.1005
R27762 VDD.n1376 VDD.n1375 1.1005
R27763 VDD.n1378 VDD.n1377 1.1005
R27764 VDD.n1318 VDD.n1317 1.1005
R27765 VDD.n1316 VDD.n1301 1.1005
R27766 VDD.n1394 VDD.n1393 1.1005
R27767 VDD.n1293 VDD.n952 1.1005
R27768 VDD.n1399 VDD.n1398 1.1005
R27769 VDD.n1292 VDD.n1291 1.1005
R27770 VDD.n1289 VDD.n952 1.1005
R27771 VDD.n1287 VDD.n1286 1.1005
R27772 VDD.n1284 VDD.n1283 1.1005
R27773 VDD.n1282 VDD.n956 1.1005
R27774 VDD.n1279 VDD.n957 1.1005
R27775 VDD.n1273 VDD.n958 1.1005
R27776 VDD.n960 VDD.n959 1.1005
R27777 VDD.n1267 VDD.n1266 1.1005
R27778 VDD.n1265 VDD.n962 1.1005
R27779 VDD.n1260 VDD.n1259 1.1005
R27780 VDD.n1249 VDD.n1248 1.1005
R27781 VDD.n1247 VDD.n967 1.1005
R27782 VDD.n1239 VDD.n968 1.1005
R27783 VDD.n1237 VDD.n1236 1.1005
R27784 VDD.n1235 VDD.n971 1.1005
R27785 VDD.n1234 VDD.n1233 1.1005
R27786 VDD.n974 VDD.n973 1.1005
R27787 VDD.n1216 VDD.n978 1.1005
R27788 VDD.n1215 VDD.n1214 1.1005
R27789 VDD.n980 VDD.n979 1.1005
R27790 VDD.n1207 VDD.n1206 1.1005
R27791 VDD.n1205 VDD.n983 1.1005
R27792 VDD.n1204 VDD.n1203 1.1005
R27793 VDD.n1201 VDD.n1200 1.1005
R27794 VDD.n1195 VDD.n985 1.1005
R27795 VDD.n1192 VDD.n986 1.1005
R27796 VDD.n1189 VDD.n987 1.1005
R27797 VDD.n1183 VDD.n988 1.1005
R27798 VDD.n1182 VDD.n1181 1.1005
R27799 VDD.n990 VDD.n989 1.1005
R27800 VDD.n1174 VDD.n1173 1.1005
R27801 VDD.n1165 VDD.n1164 1.1005
R27802 VDD.n1163 VDD.n996 1.1005
R27803 VDD.n1160 VDD.n1159 1.1005
R27804 VDD.n1156 VDD.n1155 1.1005
R27805 VDD.n1149 VDD.n1002 1.1005
R27806 VDD.n1151 VDD.n1150 1.1005
R27807 VDD.n1148 VDD.n1001 1.1005
R27808 VDD.n1140 VDD.n1007 1.1005
R27809 VDD.n1135 VDD.n1134 1.1005
R27810 VDD.n1133 VDD.n1009 1.1005
R27811 VDD.n1130 VDD.n1010 1.1005
R27812 VDD.n1124 VDD.n1123 1.1005
R27813 VDD.n1120 VDD.n1119 1.1005
R27814 VDD.n1118 VDD.n1014 1.1005
R27815 VDD.n1117 VDD.n1116 1.1005
R27816 VDD.n1017 VDD.n1016 1.1005
R27817 VDD.n1099 VDD.n1021 1.1005
R27818 VDD.n1098 VDD.n1097 1.1005
R27819 VDD.n1023 VDD.n1022 1.1005
R27820 VDD.n1090 VDD.n1089 1.1005
R27821 VDD.n1088 VDD.n1026 1.1005
R27822 VDD.n1087 VDD.n1086 1.1005
R27823 VDD.n1084 VDD.n1083 1.1005
R27824 VDD.n1078 VDD.n1028 1.1005
R27825 VDD.n1075 VDD.n1029 1.1005
R27826 VDD.n1072 VDD.n1030 1.1005
R27827 VDD.n1066 VDD.n1031 1.1005
R27828 VDD.n1065 VDD.n1064 1.1005
R27829 VDD.n1033 VDD.n1032 1.1005
R27830 VDD.n1057 VDD.n1056 1.1005
R27831 VDD.n1055 VDD.n1035 1.1005
R27832 VDD.n1049 VDD.n1036 1.1005
R27833 VDD.n1048 VDD.n1038 1.1005
R27834 VDD.n1047 VDD.n1046 1.1005
R27835 VDD.n1043 VDD.n1042 1.1005
R27836 VDD.n914 VDD.n913 1.1005
R27837 VDD.n1447 VDD.n912 1.1005
R27838 VDD.n1449 VDD.n1448 1.1005
R27839 VDD.n1450 VDD.n908 1.1005
R27840 VDD.n1455 VDD.n906 1.1005
R27841 VDD.n904 VDD.n903 1.1005
R27842 VDD.n902 VDD.n885 1.1005
R27843 VDD.n901 VDD.n900 1.1005
R27844 VDD.n1457 VDD.n1456 1.1005
R27845 VDD.n1458 VDD.n884 1.1005
R27846 VDD.n1460 VDD.n1459 1.1005
R27847 VDD.n905 VDD.n883 1.1005
R27848 VDD.n1454 VDD.n1453 1.1005
R27849 VDD.n1452 VDD.n1451 1.1005
R27850 VDD.n1446 VDD.n1445 1.1005
R27851 VDD.n1041 VDD.n1040 1.1005
R27852 VDD.n1044 VDD.n1039 1.1005
R27853 VDD.n1051 VDD.n1050 1.1005
R27854 VDD.n1058 VDD.n1034 1.1005
R27855 VDD.n1060 VDD.n1059 1.1005
R27856 VDD.n1068 VDD.n1067 1.1005
R27857 VDD.n1074 VDD.n1073 1.1005
R27858 VDD.n1077 VDD.n1076 1.1005
R27859 VDD.n1085 VDD.n1027 1.1005
R27860 VDD.n1091 VDD.n1025 1.1005
R27861 VDD.n1093 VDD.n1092 1.1005
R27862 VDD.n1101 VDD.n1100 1.1005
R27863 VDD.n1109 VDD.n1108 1.1005
R27864 VDD.n1107 VDD.n1018 1.1005
R27865 VDD.n1106 VDD.n1105 1.1005
R27866 VDD.n1020 VDD.n1019 1.1005
R27867 VDD.n1114 VDD.n1113 1.1005
R27868 VDD.n1115 VDD.n1015 1.1005
R27869 VDD.n1121 VDD.n1013 1.1005
R27870 VDD.n1122 VDD.n1011 1.1005
R27871 VDD.n1132 VDD.n1131 1.1005
R27872 VDD.n1142 VDD.n1141 1.1005
R27873 VDD.n1139 VDD.n1006 1.1005
R27874 VDD.n1138 VDD.n1137 1.1005
R27875 VDD.n1136 VDD.n1008 1.1005
R27876 VDD.n1004 VDD.n1003 1.1005
R27877 VDD.n1147 VDD.n1146 1.1005
R27878 VDD.n1000 VDD.n999 1.1005
R27879 VDD.n1157 VDD.n998 1.1005
R27880 VDD.n1158 VDD.n997 1.1005
R27881 VDD.n1172 VDD.n992 1.1005
R27882 VDD.n1167 VDD.n993 1.1005
R27883 VDD.n1169 VDD.n1168 1.1005
R27884 VDD.n1166 VDD.n995 1.1005
R27885 VDD.n1175 VDD.n991 1.1005
R27886 VDD.n1177 VDD.n1176 1.1005
R27887 VDD.n1185 VDD.n1184 1.1005
R27888 VDD.n1191 VDD.n1190 1.1005
R27889 VDD.n1194 VDD.n1193 1.1005
R27890 VDD.n1202 VDD.n984 1.1005
R27891 VDD.n1208 VDD.n982 1.1005
R27892 VDD.n1210 VDD.n1209 1.1005
R27893 VDD.n1218 VDD.n1217 1.1005
R27894 VDD.n1226 VDD.n1225 1.1005
R27895 VDD.n1224 VDD.n975 1.1005
R27896 VDD.n1223 VDD.n1222 1.1005
R27897 VDD.n977 VDD.n976 1.1005
R27898 VDD.n1231 VDD.n1230 1.1005
R27899 VDD.n1232 VDD.n972 1.1005
R27900 VDD.n1238 VDD.n970 1.1005
R27901 VDD.n1241 VDD.n1240 1.1005
R27902 VDD.n1250 VDD.n966 1.1005
R27903 VDD.n1258 VDD.n964 1.1005
R27904 VDD.n1257 VDD.n1256 1.1005
R27905 VDD.n1255 VDD.n965 1.1005
R27906 VDD.n1252 VDD.n1251 1.1005
R27907 VDD.n1261 VDD.n963 1.1005
R27908 VDD.n1264 VDD.n1263 1.1005
R27909 VDD.n1272 VDD.n1271 1.1005
R27910 VDD.n1275 VDD.n1274 1.1005
R27911 VDD.n1281 VDD.n1280 1.1005
R27912 VDD.n1291 VDD.n1290 1.1005
R27913 VDD.n1285 VDD.n955 1.1005
R27914 VDD.n1288 VDD.n951 1.1005
R27915 VDD.n893 VDD.n892 1.1005
R27916 VDD.n1473 VDD.n873 1.1005
R27917 VDD.n1498 VDD.n859 1.1005
R27918 VDD.n1555 VDD.n828 1.1005
R27919 VDD.n1581 VDD.n816 1.1005
R27920 VDD.n1606 VDD.n803 1.1005
R27921 VDD.n889 VDD.n888 1.1005
R27922 VDD.n898 VDD.n895 1.1005
R27923 VDD.n891 VDD.n874 1.1005
R27924 VDD.n1672 VDD.n771 1.1005
R27925 VDD.n1670 VDD.n1669 1.1005
R27926 VDD.n1658 VDD.n1657 1.1005
R27927 VDD.n1637 VDD.n1636 1.1005
R27928 VDD.n1633 VDD.n1632 1.1005
R27929 VDD.n1608 VDD.n1607 1.1005
R27930 VDD.n1585 VDD.n1584 1.1005
R27931 VDD.n1583 VDD.n1582 1.1005
R27932 VDD.n1559 VDD.n1558 1.1005
R27933 VDD.n1557 VDD.n1556 1.1005
R27934 VDD.n1533 VDD.n835 1.1005
R27935 VDD.n1531 VDD.n1530 1.1005
R27936 VDD.n1500 VDD.n1499 1.1005
R27937 VDD.n1477 VDD.n1476 1.1005
R27938 VDD.n1475 VDD.n1474 1.1005
R27939 VDD.n894 VDD.n887 1.1005
R27940 VDD.n896 VDD.n889 1.1005
R27941 VDD.n899 VDD.n898 1.1005
R27942 VDD.n1934 VDD.n586 1.10007
R27943 VDD.n1934 VDD.n585 1.10007
R27944 VDD.n1934 VDD.n591 1.10006
R27945 VDD.n1934 VDD.n592 1.10006
R27946 VDD.n305 VDD.n290 1.00932
R27947 VDD.n310 VDD.n283 1.00932
R27948 VDD.n299 VDD.n298 1.00926
R27949 VDD.n2026 VDD.n2019 1.00722
R27950 VDD.n2045 VDD.n2043 1.00704
R27951 VDD.n2036 VDD.n2032 1.00704
R27952 VDD.n100 VDD.n47 0.970579
R27953 VDD.n299 VDD.n297 0.941771
R27954 VDD.n310 VDD.n280 0.940947
R27955 VDD.n305 VDD.n292 0.940865
R27956 VDD.n1939 VDD.n1938 0.797844
R27957 VDD.n2045 VDD.n2023 0.738684
R27958 VDD.n1870 VDD.n673 0.733833
R27959 VDD.n1400 VDD.n1399 0.733833
R27960 VDD.n887 VDD.n886 0.733833
R27961 VDD.n1685 VDD.n765 0.733833
R27962 VDD.n460 VDD.n459 0.733833
R27963 VDD.n538 VDD.n537 0.733833
R27964 VDD.n1934 VDD.n1933 0.732782
R27965 VDD.n2042 VDD 0.668962
R27966 VDD.n2031 VDD 0.668962
R27967 VDD.n2027 VDD 0.668962
R27968 VDD.n392 VDD.n256 0.62778
R27969 VDD.n80 VDD.n79 0.62778
R27970 VDD.n806 VDD.n803 0.573769
R27971 VDD.n862 VDD.n859 0.573769
R27972 VDD.n819 VDD.n816 0.573695
R27973 VDD.n873 VDD.n871 0.573695
R27974 VDD.n831 VDD.n828 0.573346
R27975 VDD.n1561 VDD.n817 0.573297
R27976 VDD.n954 VDD.n952 0.550549
R27977 VDD.n898 VDD.n897 0.550549
R27978 VDD.n289 VDD 0.542038
R27979 VDD.n295 VDD 0.542038
R27980 VDD.n282 VDD 0.542038
R27981 VDD VDD.n253 0.533086
R27982 VDD.n1936 VDD.n576 0.4865
R27983 VDD.n253 VDD 0.41084
R27984 VDD.n1608 VDD.n802 0.39244
R27985 VDD.n1500 VDD.n858 0.39244
R27986 VDD.n1583 VDD.n815 0.389994
R27987 VDD.n1475 VDD.n872 0.389994
R27988 VDD.n1557 VDD.n827 0.387191
R27989 VDD.n1635 VDD.n787 0.384705
R27990 VDD.n1535 VDD.n1534 0.384705
R27991 VDD.n1610 VDD.n1609 0.384705
R27992 VDD.n1501 VDD.n855 0.384705
R27993 VDD.n1634 VDD.n790 0.382331
R27994 VDD.n1532 VDD.n841 0.382331
R27995 VDD.n1616 VDD.n791 0.382034
R27996 VDD.n1508 VDD.n842 0.382034
R27997 VDD.n1590 VDD.n804 0.379547
R27998 VDD.n1548 VDD.n829 0.379547
R27999 VDD.n1484 VDD.n860 0.379547
R28000 VDD.n75 VDD 0.378
R28001 VDD.n1588 VDD.n804 0.375976
R28002 VDD.n1486 VDD.n860 0.375976
R28003 VDD.n833 VDD.n829 0.375884
R28004 VDD.n1614 VDD.n791 0.374982
R28005 VDD.n1510 VDD.n842 0.374982
R28006 VDD.n1634 VDD.n788 0.374889
R28007 VDD.n1532 VDD.n840 0.374889
R28008 VDD.n1642 VDD.n1635 0.373984
R28009 VDD.n1534 VDD.n837 0.373984
R28010 VDD.n1609 VDD.n801 0.373891
R28011 VDD.n1502 VDD.n1501 0.373891
R28012 VDD.n2040 VDD.n2023 0.361965
R28013 VDD VDD.n76 0.36028
R28014 VDD.n255 VDD.n252 0.329931
R28015 VDD.n78 VDD.n71 0.329931
R28016 VDD VDD.n254 0.315825
R28017 VDD VDD.n77 0.315825
R28018 VDD.n1937 VDD.n1936 0.290686
R28019 VDD.n1565 VDD.n817 0.280767
R28020 VDD.n1673 VDD.n765 0.275034
R28021 VDD.n256 VDD 0.239511
R28022 VDD.n79 VDD 0.239511
R28023 VDD.n289 VDD.n288 0.237776
R28024 VDD.n300 VDD.n295 0.237776
R28025 VDD.n282 VDD.n281 0.237776
R28026 VDD VDD.n2030 0.236427
R28027 VDD.n2024 VDD 0.23614
R28028 VDD VDD.n2052 0.227409
R28029 VDD.n76 VDD.n75 0.222011
R28030 VDD.n2051 VDD 0.2205
R28031 VDD.n2029 VDD.n2024 0.21461
R28032 VDD.n2038 VDD.n2030 0.214316
R28033 VDD.n303 VDD.n288 0.21301
R28034 VDD.n301 VDD.n300 0.21301
R28035 VDD.n293 VDD.n281 0.21301
R28036 VDD.n297 VDD 0.211907
R28037 VDD.n292 VDD 0.21003
R28038 VDD VDD.n280 0.209914
R28039 VDD.n558 VDD.n555 0.205151
R28040 VDD.n558 VDD.n553 0.205151
R28041 VDD.n563 VDD.n553 0.205151
R28042 VDD.n557 VDD.n552 0.205151
R28043 VDD.n564 VDD.n552 0.205151
R28044 VDD.n565 VDD.n551 0.205151
R28045 VDD.n559 VDD.n554 0.202799
R28046 VDD.n311 VDD.n279 0.189575
R28047 VDD VDD.n280 0.184885
R28048 VDD VDD.n292 0.184754
R28049 VDD.n439 VDD.n435 0.183833
R28050 VDD.n447 VDD.n435 0.183833
R28051 VDD.n448 VDD.n447 0.183833
R28052 VDD.n449 VDD.n448 0.183833
R28053 VDD.n449 VDD.n427 0.183833
R28054 VDD.n459 VDD.n427 0.183833
R28055 VDD.n461 VDD.n460 0.183833
R28056 VDD.n461 VDD.n419 0.183833
R28057 VDD.n471 VDD.n419 0.183833
R28058 VDD.n472 VDD.n471 0.183833
R28059 VDD.n474 VDD.n472 0.183833
R28060 VDD.n474 VDD.n473 0.183833
R28061 VDD.n473 VDD.n410 0.183833
R28062 VDD.n485 VDD.n410 0.183833
R28063 VDD.n486 VDD.n485 0.183833
R28064 VDD.n487 VDD.n486 0.183833
R28065 VDD.n487 VDD.n408 0.183833
R28066 VDD.n492 VDD.n408 0.183833
R28067 VDD.n493 VDD.n492 0.183833
R28068 VDD.n539 VDD.n493 0.183833
R28069 VDD.n539 VDD.n538 0.183833
R28070 VDD.n537 VDD.n494 0.183833
R28071 VDD.n533 VDD.n494 0.183833
R28072 VDD.n533 VDD.n532 0.183833
R28073 VDD.n532 VDD.n531 0.183833
R28074 VDD.n531 VDD.n499 0.183833
R28075 VDD.n527 VDD.n499 0.183833
R28076 VDD.n527 VDD.n526 0.183833
R28077 VDD.n297 VDD 0.182972
R28078 VDD.n254 VDD 0.180486
R28079 VDD.n77 VDD 0.180486
R28080 VDD.n2026 VDD 0.179399
R28081 VDD VDD.n2043 0.179186
R28082 VDD VDD.n2032 0.179186
R28083 VDD.n298 VDD 0.174803
R28084 VDD.n290 VDD 0.173911
R28085 VDD.n283 VDD 0.173911
R28086 VDD.n2043 VDD.n2042 0.173371
R28087 VDD.n2032 VDD.n2031 0.173371
R28088 VDD.n2027 VDD.n2026 0.173186
R28089 VDD.n298 VDD.n295 0.17126
R28090 VDD.n290 VDD.n289 0.171175
R28091 VDD.n283 VDD.n282 0.171175
R28092 VDD.n309 VDD.n279 0.160581
R28093 VDD.n464 VDD.n424 0.149653
R28094 VDD.n464 VDD.n422 0.149653
R28095 VDD.n468 VDD.n422 0.149653
R28096 VDD.n468 VDD.n415 0.149653
R28097 VDD.n477 VDD.n415 0.149653
R28098 VDD.n477 VDD.n413 0.149653
R28099 VDD.n481 VDD.n413 0.149653
R28100 VDD.n481 VDD.n397 0.149653
R28101 VDD.n549 VDD.n397 0.149653
R28102 VDD.n549 VDD.n548 0.149653
R28103 VDD.n548 VDD.n547 0.149653
R28104 VDD.n547 VDD.n401 0.149653
R28105 VDD.n543 VDD.n401 0.149653
R28106 VDD.n543 VDD.n542 0.149653
R28107 VDD.n542 VDD.n404 0.149653
R28108 VDD.n463 VDD.n425 0.149653
R28109 VDD.n463 VDD.n421 0.149653
R28110 VDD.n469 VDD.n421 0.149653
R28111 VDD.n469 VDD.n416 0.149653
R28112 VDD.n476 VDD.n416 0.149653
R28113 VDD.n476 VDD.n412 0.149653
R28114 VDD.n482 VDD.n412 0.149653
R28115 VDD.n483 VDD.n482 0.149653
R28116 VDD.n483 VDD.n398 0.149653
R28117 VDD.n399 VDD.n398 0.149653
R28118 VDD.n400 VDD.n399 0.149653
R28119 VDD.n490 VDD.n400 0.149653
R28120 VDD.n490 VDD.n403 0.149653
R28121 VDD.n541 VDD.n403 0.149653
R28122 VDD.n541 VDD.n405 0.149653
R28123 VDD.n462 VDD.n426 0.149653
R28124 VDD.n462 VDD.n420 0.149653
R28125 VDD.n470 VDD.n420 0.149653
R28126 VDD.n470 VDD.n417 0.149653
R28127 VDD.n475 VDD.n417 0.149653
R28128 VDD.n475 VDD.n418 0.149653
R28129 VDD.n418 VDD.n411 0.149653
R28130 VDD.n484 VDD.n411 0.149653
R28131 VDD.n484 VDD.n409 0.149653
R28132 VDD.n488 VDD.n409 0.149653
R28133 VDD.n489 VDD.n488 0.149653
R28134 VDD.n491 VDD.n489 0.149653
R28135 VDD.n491 VDD.n406 0.149653
R28136 VDD.n540 VDD.n406 0.149653
R28137 VDD.n540 VDD.n407 0.149653
R28138 VDD.n440 VDD.n436 0.149653
R28139 VDD.n446 VDD.n436 0.149653
R28140 VDD.n446 VDD.n434 0.149653
R28141 VDD.n450 VDD.n434 0.149653
R28142 VDD.n450 VDD.n428 0.149653
R28143 VDD.n458 VDD.n428 0.149653
R28144 VDD.n441 VDD.n437 0.149653
R28145 VDD.n445 VDD.n437 0.149653
R28146 VDD.n445 VDD.n433 0.149653
R28147 VDD.n451 VDD.n433 0.149653
R28148 VDD.n451 VDD.n429 0.149653
R28149 VDD.n457 VDD.n429 0.149653
R28150 VDD.n444 VDD.n438 0.149653
R28151 VDD.n444 VDD.n432 0.149653
R28152 VDD.n452 VDD.n432 0.149653
R28153 VDD.n452 VDD.n430 0.149653
R28154 VDD.n456 VDD.n430 0.149653
R28155 VDD.n526 VDD.n525 0.149
R28156 VDD.n513 VDD.n512 0.147167
R28157 VDD.n514 VDD.n513 0.147167
R28158 VDD.n514 VDD.n508 0.147167
R28159 VDD.n518 VDD.n508 0.147167
R28160 VDD.n519 VDD.n518 0.147167
R28161 VDD.n520 VDD.n519 0.147167
R28162 VDD.n520 VDD.n505 0.147167
R28163 VDD.n496 VDD.n495 0.147167
R28164 VDD.n497 VDD.n496 0.147167
R28165 VDD.n507 VDD.n497 0.147167
R28166 VDD.n507 VDD.n500 0.147167
R28167 VDD.n501 VDD.n500 0.147167
R28168 VDD.n502 VDD.n501 0.147167
R28169 VDD.n504 VDD.n502 0.147167
R28170 VDD.n523 VDD.n504 0.147167
R28171 VDD.n536 VDD.n535 0.147167
R28172 VDD.n535 VDD.n534 0.147167
R28173 VDD.n534 VDD.n498 0.147167
R28174 VDD.n530 VDD.n498 0.147167
R28175 VDD.n530 VDD.n529 0.147167
R28176 VDD.n529 VDD.n528 0.147167
R28177 VDD.n528 VDD.n503 0.147167
R28178 VDD.n524 VDD.n503 0.147167
R28179 VDD.n2052 VDD.n2051 0.142085
R28180 VDD.n314 VDD.n313 0.138
R28181 VDD.n315 VDD.n314 0.138
R28182 VDD.n315 VDD.n277 0.138
R28183 VDD.n320 VDD.n277 0.138
R28184 VDD.n321 VDD.n320 0.138
R28185 VDD.n322 VDD.n321 0.138
R28186 VDD.n322 VDD.n275 0.138
R28187 VDD.n327 VDD.n275 0.138
R28188 VDD.n328 VDD.n327 0.138
R28189 VDD.n329 VDD.n328 0.138
R28190 VDD.n329 VDD.n273 0.138
R28191 VDD.n334 VDD.n273 0.138
R28192 VDD.n335 VDD.n334 0.138
R28193 VDD.n336 VDD.n335 0.138
R28194 VDD.n336 VDD.n271 0.138
R28195 VDD.n341 VDD.n271 0.138
R28196 VDD.n342 VDD.n341 0.138
R28197 VDD.n343 VDD.n342 0.138
R28198 VDD.n343 VDD.n269 0.138
R28199 VDD.n348 VDD.n269 0.138
R28200 VDD.n349 VDD.n348 0.138
R28201 VDD.n350 VDD.n349 0.138
R28202 VDD.n350 VDD.n267 0.138
R28203 VDD.n355 VDD.n267 0.138
R28204 VDD.n356 VDD.n355 0.138
R28205 VDD.n357 VDD.n356 0.138
R28206 VDD.n357 VDD.n265 0.138
R28207 VDD.n362 VDD.n265 0.138
R28208 VDD.n363 VDD.n362 0.138
R28209 VDD.n364 VDD.n363 0.138
R28210 VDD.n364 VDD.n263 0.138
R28211 VDD.n369 VDD.n263 0.138
R28212 VDD.n370 VDD.n369 0.138
R28213 VDD.n371 VDD.n370 0.138
R28214 VDD.n371 VDD.n261 0.138
R28215 VDD.n376 VDD.n261 0.138
R28216 VDD.n377 VDD.n376 0.138
R28217 VDD.n378 VDD.n377 0.138
R28218 VDD.n378 VDD.n259 0.138
R28219 VDD.n383 VDD.n259 0.138
R28220 VDD.n384 VDD.n383 0.138
R28221 VDD.n385 VDD.n384 0.138
R28222 VDD.n385 VDD.n257 0.138
R28223 VDD.n390 VDD.n257 0.138
R28224 VDD.n391 VDD.n390 0.138
R28225 VDD.n81 VDD.n65 0.138
R28226 VDD.n91 VDD.n65 0.138
R28227 VDD.n92 VDD.n91 0.138
R28228 VDD.n94 VDD.n92 0.138
R28229 VDD.n94 VDD.n93 0.138
R28230 VDD.n93 VDD.n57 0.138
R28231 VDD.n105 VDD.n57 0.138
R28232 VDD.n106 VDD.n105 0.138
R28233 VDD.n107 VDD.n106 0.138
R28234 VDD.n107 VDD.n55 0.138
R28235 VDD.n111 VDD.n55 0.138
R28236 VDD.n112 VDD.n111 0.138
R28237 VDD.n113 VDD.n112 0.138
R28238 VDD.n113 VDD.n53 0.138
R28239 VDD.n117 VDD.n53 0.138
R28240 VDD.n118 VDD.n117 0.138
R28241 VDD.n119 VDD.n118 0.138
R28242 VDD.n119 VDD.n51 0.138
R28243 VDD.n123 VDD.n51 0.138
R28244 VDD.n124 VDD.n123 0.138
R28245 VDD.n125 VDD.n124 0.138
R28246 VDD.n125 VDD.n43 0.138
R28247 VDD.n135 VDD.n43 0.138
R28248 VDD.n136 VDD.n135 0.138
R28249 VDD.n137 VDD.n136 0.138
R28250 VDD.n137 VDD.n35 0.138
R28251 VDD.n147 VDD.n35 0.138
R28252 VDD.n148 VDD.n147 0.138
R28253 VDD.n149 VDD.n148 0.138
R28254 VDD.n149 VDD.n27 0.138
R28255 VDD.n159 VDD.n27 0.138
R28256 VDD.n160 VDD.n159 0.138
R28257 VDD.n161 VDD.n160 0.138
R28258 VDD.n161 VDD.n19 0.138
R28259 VDD.n171 VDD.n19 0.138
R28260 VDD.n172 VDD.n171 0.138
R28261 VDD.n173 VDD.n172 0.138
R28262 VDD.n173 VDD.n11 0.138
R28263 VDD.n184 VDD.n11 0.138
R28264 VDD.n185 VDD.n184 0.138
R28265 VDD.n186 VDD.n185 0.138
R28266 VDD.n186 VDD.n2 0.138
R28267 VDD.n2017 VDD.n2 0.138
R28268 VDD.n2018 VDD.n2017 0.138
R28269 VDD.n2053 VDD.n2018 0.138
R28270 VDD.n1938 VDD.n1937 0.125553
R28271 VDD.n72 VDD 0.120789
R28272 VDD.n439 VDD 0.114167
R28273 VDD.n392 VDD.n391 0.11325
R28274 VDD.n81 VDD.n80 0.11325
R28275 VDD.n195 VDD.n194 0.111892
R28276 VDD.n196 VDD.n195 0.111892
R28277 VDD.n317 VDD.n196 0.111892
R28278 VDD.n317 VDD.n199 0.111892
R28279 VDD.n200 VDD.n199 0.111892
R28280 VDD.n201 VDD.n200 0.111892
R28281 VDD.n324 VDD.n201 0.111892
R28282 VDD.n324 VDD.n204 0.111892
R28283 VDD.n205 VDD.n204 0.111892
R28284 VDD.n206 VDD.n205 0.111892
R28285 VDD.n331 VDD.n206 0.111892
R28286 VDD.n331 VDD.n209 0.111892
R28287 VDD.n210 VDD.n209 0.111892
R28288 VDD.n211 VDD.n210 0.111892
R28289 VDD.n338 VDD.n211 0.111892
R28290 VDD.n338 VDD.n214 0.111892
R28291 VDD.n215 VDD.n214 0.111892
R28292 VDD.n216 VDD.n215 0.111892
R28293 VDD.n345 VDD.n216 0.111892
R28294 VDD.n345 VDD.n219 0.111892
R28295 VDD.n220 VDD.n219 0.111892
R28296 VDD.n221 VDD.n220 0.111892
R28297 VDD.n352 VDD.n221 0.111892
R28298 VDD.n352 VDD.n224 0.111892
R28299 VDD.n225 VDD.n224 0.111892
R28300 VDD.n226 VDD.n225 0.111892
R28301 VDD.n359 VDD.n226 0.111892
R28302 VDD.n359 VDD.n229 0.111892
R28303 VDD.n230 VDD.n229 0.111892
R28304 VDD.n231 VDD.n230 0.111892
R28305 VDD.n366 VDD.n231 0.111892
R28306 VDD.n366 VDD.n234 0.111892
R28307 VDD.n235 VDD.n234 0.111892
R28308 VDD.n236 VDD.n235 0.111892
R28309 VDD.n373 VDD.n236 0.111892
R28310 VDD.n373 VDD.n239 0.111892
R28311 VDD.n240 VDD.n239 0.111892
R28312 VDD.n241 VDD.n240 0.111892
R28313 VDD.n380 VDD.n241 0.111892
R28314 VDD.n380 VDD.n244 0.111892
R28315 VDD.n245 VDD.n244 0.111892
R28316 VDD.n246 VDD.n245 0.111892
R28317 VDD.n387 VDD.n246 0.111892
R28318 VDD.n387 VDD.n249 0.111892
R28319 VDD.n250 VDD.n249 0.111892
R28320 VDD.n394 VDD.n250 0.111892
R28321 VDD.n2009 VDD.n2008 0.111892
R28322 VDD.n2008 VDD.n2007 0.111892
R28323 VDD.n2007 VDD.n197 0.111892
R28324 VDD.n2003 VDD.n197 0.111892
R28325 VDD.n2003 VDD.n2002 0.111892
R28326 VDD.n2002 VDD.n2001 0.111892
R28327 VDD.n2001 VDD.n202 0.111892
R28328 VDD.n1997 VDD.n202 0.111892
R28329 VDD.n1997 VDD.n1996 0.111892
R28330 VDD.n1996 VDD.n1995 0.111892
R28331 VDD.n1995 VDD.n207 0.111892
R28332 VDD.n1991 VDD.n207 0.111892
R28333 VDD.n1991 VDD.n1990 0.111892
R28334 VDD.n1990 VDD.n1989 0.111892
R28335 VDD.n1989 VDD.n212 0.111892
R28336 VDD.n1985 VDD.n212 0.111892
R28337 VDD.n1985 VDD.n1984 0.111892
R28338 VDD.n1984 VDD.n1983 0.111892
R28339 VDD.n1983 VDD.n217 0.111892
R28340 VDD.n1979 VDD.n217 0.111892
R28341 VDD.n1979 VDD.n1978 0.111892
R28342 VDD.n1978 VDD.n1977 0.111892
R28343 VDD.n1977 VDD.n222 0.111892
R28344 VDD.n1973 VDD.n222 0.111892
R28345 VDD.n1973 VDD.n1972 0.111892
R28346 VDD.n1972 VDD.n1971 0.111892
R28347 VDD.n1971 VDD.n227 0.111892
R28348 VDD.n1967 VDD.n227 0.111892
R28349 VDD.n1967 VDD.n1966 0.111892
R28350 VDD.n1966 VDD.n1965 0.111892
R28351 VDD.n1965 VDD.n232 0.111892
R28352 VDD.n1961 VDD.n232 0.111892
R28353 VDD.n1961 VDD.n1960 0.111892
R28354 VDD.n1960 VDD.n1959 0.111892
R28355 VDD.n1959 VDD.n237 0.111892
R28356 VDD.n1955 VDD.n237 0.111892
R28357 VDD.n1955 VDD.n1954 0.111892
R28358 VDD.n1954 VDD.n1953 0.111892
R28359 VDD.n1953 VDD.n242 0.111892
R28360 VDD.n1949 VDD.n242 0.111892
R28361 VDD.n1949 VDD.n1948 0.111892
R28362 VDD.n1948 VDD.n1947 0.111892
R28363 VDD.n1947 VDD.n247 0.111892
R28364 VDD.n1943 VDD.n247 0.111892
R28365 VDD.n1943 VDD.n1942 0.111892
R28366 VDD.n1942 VDD.n1941 0.111892
R28367 VDD.n279 VDD 0.11175
R28368 VDD.n312 VDD.n278 0.1105
R28369 VDD.n316 VDD.n278 0.1105
R28370 VDD.n318 VDD.n316 0.1105
R28371 VDD.n319 VDD.n318 0.1105
R28372 VDD.n319 VDD.n276 0.1105
R28373 VDD.n323 VDD.n276 0.1105
R28374 VDD.n325 VDD.n323 0.1105
R28375 VDD.n326 VDD.n325 0.1105
R28376 VDD.n326 VDD.n274 0.1105
R28377 VDD.n330 VDD.n274 0.1105
R28378 VDD.n332 VDD.n330 0.1105
R28379 VDD.n333 VDD.n332 0.1105
R28380 VDD.n333 VDD.n272 0.1105
R28381 VDD.n337 VDD.n272 0.1105
R28382 VDD.n339 VDD.n337 0.1105
R28383 VDD.n340 VDD.n339 0.1105
R28384 VDD.n340 VDD.n270 0.1105
R28385 VDD.n344 VDD.n270 0.1105
R28386 VDD.n346 VDD.n344 0.1105
R28387 VDD.n347 VDD.n346 0.1105
R28388 VDD.n347 VDD.n268 0.1105
R28389 VDD.n351 VDD.n268 0.1105
R28390 VDD.n353 VDD.n351 0.1105
R28391 VDD.n354 VDD.n353 0.1105
R28392 VDD.n354 VDD.n266 0.1105
R28393 VDD.n358 VDD.n266 0.1105
R28394 VDD.n360 VDD.n358 0.1105
R28395 VDD.n361 VDD.n360 0.1105
R28396 VDD.n361 VDD.n264 0.1105
R28397 VDD.n365 VDD.n264 0.1105
R28398 VDD.n367 VDD.n365 0.1105
R28399 VDD.n368 VDD.n367 0.1105
R28400 VDD.n368 VDD.n262 0.1105
R28401 VDD.n372 VDD.n262 0.1105
R28402 VDD.n374 VDD.n372 0.1105
R28403 VDD.n375 VDD.n374 0.1105
R28404 VDD.n375 VDD.n260 0.1105
R28405 VDD.n379 VDD.n260 0.1105
R28406 VDD.n381 VDD.n379 0.1105
R28407 VDD.n382 VDD.n381 0.1105
R28408 VDD.n382 VDD.n258 0.1105
R28409 VDD.n386 VDD.n258 0.1105
R28410 VDD.n388 VDD.n386 0.1105
R28411 VDD.n389 VDD.n388 0.1105
R28412 VDD.n389 VDD.n251 0.1105
R28413 VDD.n393 VDD.n251 0.1105
R28414 VDD.n128 VDD.n48 0.1105
R28415 VDD.n128 VDD.n46 0.1105
R28416 VDD.n132 VDD.n46 0.1105
R28417 VDD.n132 VDD.n40 0.1105
R28418 VDD.n140 VDD.n40 0.1105
R28419 VDD.n140 VDD.n38 0.1105
R28420 VDD.n144 VDD.n38 0.1105
R28421 VDD.n144 VDD.n32 0.1105
R28422 VDD.n152 VDD.n32 0.1105
R28423 VDD.n152 VDD.n30 0.1105
R28424 VDD.n156 VDD.n30 0.1105
R28425 VDD.n156 VDD.n24 0.1105
R28426 VDD.n164 VDD.n24 0.1105
R28427 VDD.n164 VDD.n22 0.1105
R28428 VDD.n168 VDD.n22 0.1105
R28429 VDD.n168 VDD.n16 0.1105
R28430 VDD.n176 VDD.n16 0.1105
R28431 VDD.n176 VDD.n14 0.1105
R28432 VDD.n181 VDD.n14 0.1105
R28433 VDD.n181 VDD.n8 0.1105
R28434 VDD.n189 VDD.n8 0.1105
R28435 VDD.n190 VDD.n189 0.1105
R28436 VDD.n190 VDD.n5 0.1105
R28437 VDD.n2013 VDD.n5 0.1105
R28438 VDD.n2013 VDD.n6 0.1105
R28439 VDD.n127 VDD.n49 0.1105
R28440 VDD.n127 VDD.n45 0.1105
R28441 VDD.n133 VDD.n45 0.1105
R28442 VDD.n133 VDD.n41 0.1105
R28443 VDD.n139 VDD.n41 0.1105
R28444 VDD.n139 VDD.n37 0.1105
R28445 VDD.n145 VDD.n37 0.1105
R28446 VDD.n145 VDD.n33 0.1105
R28447 VDD.n151 VDD.n33 0.1105
R28448 VDD.n151 VDD.n29 0.1105
R28449 VDD.n157 VDD.n29 0.1105
R28450 VDD.n157 VDD.n25 0.1105
R28451 VDD.n163 VDD.n25 0.1105
R28452 VDD.n163 VDD.n21 0.1105
R28453 VDD.n169 VDD.n21 0.1105
R28454 VDD.n169 VDD.n17 0.1105
R28455 VDD.n175 VDD.n17 0.1105
R28456 VDD.n175 VDD.n13 0.1105
R28457 VDD.n182 VDD.n13 0.1105
R28458 VDD.n182 VDD.n9 0.1105
R28459 VDD.n188 VDD.n9 0.1105
R28460 VDD.n188 VDD.n4 0.1105
R28461 VDD.n2015 VDD.n4 0.1105
R28462 VDD.n2015 VDD.n2014 0.1105
R28463 VDD.n2014 VDD.n1 0.1105
R28464 VDD.n82 VDD.n70 0.1105
R28465 VDD.n82 VDD.n66 0.1105
R28466 VDD.n90 VDD.n66 0.1105
R28467 VDD.n90 VDD.n64 0.1105
R28468 VDD.n95 VDD.n64 0.1105
R28469 VDD.n95 VDD.n58 0.1105
R28470 VDD.n103 VDD.n58 0.1105
R28471 VDD.n104 VDD.n103 0.1105
R28472 VDD.n104 VDD.n56 0.1105
R28473 VDD.n108 VDD.n56 0.1105
R28474 VDD.n109 VDD.n108 0.1105
R28475 VDD.n110 VDD.n109 0.1105
R28476 VDD.n110 VDD.n54 0.1105
R28477 VDD.n114 VDD.n54 0.1105
R28478 VDD.n115 VDD.n114 0.1105
R28479 VDD.n116 VDD.n115 0.1105
R28480 VDD.n116 VDD.n52 0.1105
R28481 VDD.n120 VDD.n52 0.1105
R28482 VDD.n121 VDD.n120 0.1105
R28483 VDD.n122 VDD.n121 0.1105
R28484 VDD.n122 VDD.n50 0.1105
R28485 VDD.n126 VDD.n50 0.1105
R28486 VDD.n126 VDD.n44 0.1105
R28487 VDD.n134 VDD.n44 0.1105
R28488 VDD.n134 VDD.n42 0.1105
R28489 VDD.n138 VDD.n42 0.1105
R28490 VDD.n138 VDD.n36 0.1105
R28491 VDD.n146 VDD.n36 0.1105
R28492 VDD.n146 VDD.n34 0.1105
R28493 VDD.n150 VDD.n34 0.1105
R28494 VDD.n150 VDD.n28 0.1105
R28495 VDD.n158 VDD.n28 0.1105
R28496 VDD.n158 VDD.n26 0.1105
R28497 VDD.n162 VDD.n26 0.1105
R28498 VDD.n162 VDD.n20 0.1105
R28499 VDD.n170 VDD.n20 0.1105
R28500 VDD.n170 VDD.n18 0.1105
R28501 VDD.n174 VDD.n18 0.1105
R28502 VDD.n174 VDD.n12 0.1105
R28503 VDD.n183 VDD.n12 0.1105
R28504 VDD.n183 VDD.n10 0.1105
R28505 VDD.n187 VDD.n10 0.1105
R28506 VDD.n187 VDD.n3 0.1105
R28507 VDD.n2016 VDD.n3 0.1105
R28508 VDD.n2016 VDD.n0 0.1105
R28509 VDD.n2054 VDD.n0 0.1105
R28510 VDD.n84 VDD.n83 0.1105
R28511 VDD.n83 VDD.n67 0.1105
R28512 VDD.n89 VDD.n67 0.1105
R28513 VDD.n89 VDD.n63 0.1105
R28514 VDD.n96 VDD.n63 0.1105
R28515 VDD.n96 VDD.n59 0.1105
R28516 VDD.n102 VDD.n59 0.1105
R28517 VDD.n69 VDD.n68 0.1105
R28518 VDD.n88 VDD.n68 0.1105
R28519 VDD.n88 VDD.n62 0.1105
R28520 VDD.n97 VDD.n62 0.1105
R28521 VDD.n97 VDD.n60 0.1105
R28522 VDD.n101 VDD.n60 0.1105
R28523 VDD.n73 VDD.n72 0.108289
R28524 VDD.n562 VDD.n561 0.102356
R28525 VDD.n557 VDD.n556 0.101051
R28526 VDD.n561 VDD.n554 0.0997237
R28527 VDD.n560 VDD.n559 0.0997007
R28528 VDD.n571 VDD.n568 0.0965
R28529 VDD.n573 VDD.n567 0.0965
R28530 VDD.n573 VDD.n572 0.0965
R28531 VDD.n575 VDD.n574 0.0965
R28532 VDD.n309 VDD.n308 0.0929625
R28533 VDD.n1936 VDD.n1935 0.0806174
R28534 VDD VDD.n2022 0.0805073
R28535 VDD VDD.n2033 0.0805073
R28536 VDD VDD.n2020 0.0805073
R28537 VDD.n1935 VDD 0.0792814
R28538 VDD.n393 VDD 0.0775
R28539 VDD VDD.n2054 0.0775
R28540 VDD.n2023 VDD 0.075162
R28541 VDD.n442 VDD.n438 0.0749488
R28542 VDD.n522 VDD.n505 0.0737263
R28543 VDD.n87 VDD.n86 0.0697913
R28544 VDD.n87 VDD.n61 0.0697913
R28545 VDD.n98 VDD.n61 0.0697913
R28546 VDD.n99 VDD.n98 0.0697913
R28547 VDD.n100 VDD.n99 0.0697913
R28548 VDD.n129 VDD.n47 0.0697913
R28549 VDD.n130 VDD.n129 0.0697913
R28550 VDD.n131 VDD.n130 0.0697913
R28551 VDD.n131 VDD.n39 0.0697913
R28552 VDD.n141 VDD.n39 0.0697913
R28553 VDD.n142 VDD.n141 0.0697913
R28554 VDD.n143 VDD.n142 0.0697913
R28555 VDD.n143 VDD.n31 0.0697913
R28556 VDD.n153 VDD.n31 0.0697913
R28557 VDD.n154 VDD.n153 0.0697913
R28558 VDD.n155 VDD.n154 0.0697913
R28559 VDD.n155 VDD.n23 0.0697913
R28560 VDD.n165 VDD.n23 0.0697913
R28561 VDD.n166 VDD.n165 0.0697913
R28562 VDD.n167 VDD.n166 0.0697913
R28563 VDD.n167 VDD.n15 0.0697913
R28564 VDD.n177 VDD.n15 0.0697913
R28565 VDD.n178 VDD.n177 0.0697913
R28566 VDD.n180 VDD.n178 0.0697913
R28567 VDD.n180 VDD.n179 0.0697913
R28568 VDD.n179 VDD.n7 0.0697913
R28569 VDD.n191 VDD.n7 0.0697913
R28570 VDD.n192 VDD.n191 0.0697913
R28571 VDD.n2012 VDD.n192 0.0697913
R28572 VDD.n2012 VDD.n2011 0.0697913
R28573 VDD.n2010 VDD.n193 0.0697913
R28574 VDD.n2006 VDD.n193 0.0697913
R28575 VDD.n2006 VDD.n2005 0.0697913
R28576 VDD.n2005 VDD.n2004 0.0697913
R28577 VDD.n2004 VDD.n198 0.0697913
R28578 VDD.n2000 VDD.n198 0.0697913
R28579 VDD.n2000 VDD.n1999 0.0697913
R28580 VDD.n1999 VDD.n1998 0.0697913
R28581 VDD.n1998 VDD.n203 0.0697913
R28582 VDD.n1994 VDD.n203 0.0697913
R28583 VDD.n1994 VDD.n1993 0.0697913
R28584 VDD.n1993 VDD.n1992 0.0697913
R28585 VDD.n1992 VDD.n208 0.0697913
R28586 VDD.n1988 VDD.n208 0.0697913
R28587 VDD.n1988 VDD.n1987 0.0697913
R28588 VDD.n1987 VDD.n1986 0.0697913
R28589 VDD.n1986 VDD.n213 0.0697913
R28590 VDD.n1982 VDD.n213 0.0697913
R28591 VDD.n1982 VDD.n1981 0.0697913
R28592 VDD.n1981 VDD.n1980 0.0697913
R28593 VDD.n1980 VDD.n218 0.0697913
R28594 VDD.n1976 VDD.n218 0.0697913
R28595 VDD.n1976 VDD.n1975 0.0697913
R28596 VDD.n1975 VDD.n1974 0.0697913
R28597 VDD.n1974 VDD.n223 0.0697913
R28598 VDD.n1970 VDD.n223 0.0697913
R28599 VDD.n1970 VDD.n1969 0.0697913
R28600 VDD.n1969 VDD.n1968 0.0697913
R28601 VDD.n1968 VDD.n228 0.0697913
R28602 VDD.n1964 VDD.n228 0.0697913
R28603 VDD.n1964 VDD.n1963 0.0697913
R28604 VDD.n1963 VDD.n1962 0.0697913
R28605 VDD.n1962 VDD.n233 0.0697913
R28606 VDD.n1958 VDD.n233 0.0697913
R28607 VDD.n1958 VDD.n1957 0.0697913
R28608 VDD.n1957 VDD.n1956 0.0697913
R28609 VDD.n1956 VDD.n238 0.0697913
R28610 VDD.n1952 VDD.n238 0.0697913
R28611 VDD.n1952 VDD.n1951 0.0697913
R28612 VDD.n1951 VDD.n1950 0.0697913
R28613 VDD.n1950 VDD.n243 0.0697913
R28614 VDD.n1946 VDD.n243 0.0697913
R28615 VDD.n1946 VDD.n1945 0.0697913
R28616 VDD.n1945 VDD.n1944 0.0697913
R28617 VDD.n1944 VDD.n248 0.0697913
R28618 VDD.n1940 VDD.n248 0.0697913
R28619 VDD.n2047 VDD.n2022 0.0668943
R28620 VDD.n2033 VDD.n2021 0.0668943
R28621 VDD.n2049 VDD.n2020 0.0668943
R28622 VDD.n73 VDD 0.0661393
R28623 VDD VDD.n287 0.0623351
R28624 VDD.n306 VDD 0.0619977
R28625 VDD.n570 VDD 0.0605
R28626 VDD.n304 VDD.n303 0.0569103
R28627 VDD.n301 VDD.n294 0.0569103
R28628 VDD.n293 VDD.n284 0.0569103
R28629 VDD.n2041 VDD.n2040 0.0569103
R28630 VDD.n2038 VDD.n2037 0.0569103
R28631 VDD.n2029 VDD.n2028 0.0569103
R28632 VDD.n85 VDD.n69 0.0554576
R28633 VDD.n279 VDD 0.054882
R28634 VDD.n2051 VDD 0.054882
R28635 VDD VDD.n285 0.0539078
R28636 VDD.n308 VDD.n286 0.053691
R28637 VDD.n291 VDD 0.0535728
R28638 VDD.n296 VDD 0.0535728
R28639 VDD VDD.n1934 0.0506457
R28640 VDD.n525 VDD 0.05
R28641 VDD VDD.n2025 0.0484979
R28642 VDD.n574 VDD.n566 0.0484934
R28643 VDD.n569 VDD.n568 0.0484338
R28644 VDD.n2044 VDD 0.0481629
R28645 VDD.n2035 VDD 0.0481629
R28646 VDD.n286 VDD 0.0442237
R28647 VDD.n304 VDD 0.0428077
R28648 VDD VDD.n294 0.0428077
R28649 VDD.n284 VDD 0.0428077
R28650 VDD.n2042 VDD.n2041 0.0428077
R28651 VDD.n2037 VDD.n2031 0.0428077
R28652 VDD.n2028 VDD.n2027 0.0428077
R28653 VDD.n1463 VDD.n880 0.0405
R28654 VDD.n1441 VDD.n880 0.0405
R28655 VDD.n1441 VDD.n916 0.0405
R28656 VDD.n1437 VDD.n916 0.0405
R28657 VDD.n1437 VDD.n1436 0.0405
R28658 VDD.n1436 VDD.n1435 0.0405
R28659 VDD.n1435 VDD.n921 0.0405
R28660 VDD.n1431 VDD.n921 0.0405
R28661 VDD.n1431 VDD.n1430 0.0405
R28662 VDD.n1430 VDD.n1429 0.0405
R28663 VDD.n1429 VDD.n926 0.0405
R28664 VDD.n1425 VDD.n926 0.0405
R28665 VDD.n1425 VDD.n1424 0.0405
R28666 VDD.n1424 VDD.n1423 0.0405
R28667 VDD.n1419 VDD.n931 0.0405
R28668 VDD.n1419 VDD.n1418 0.0405
R28669 VDD.n1418 VDD.n1417 0.0405
R28670 VDD.n1417 VDD.n936 0.0405
R28671 VDD.n1413 VDD.n936 0.0405
R28672 VDD.n1413 VDD.n1412 0.0405
R28673 VDD.n1412 VDD.n1411 0.0405
R28674 VDD.n1411 VDD.n941 0.0405
R28675 VDD.n1407 VDD.n941 0.0405
R28676 VDD.n1407 VDD.n1406 0.0405
R28677 VDD.n1406 VDD.n1405 0.0405
R28678 VDD.n1405 VDD.n946 0.0405
R28679 VDD.n1699 VDD.n749 0.0405
R28680 VDD.n1700 VDD.n1699 0.0405
R28681 VDD.n1701 VDD.n1700 0.0405
R28682 VDD.n1701 VDD.n737 0.0405
R28683 VDD.n1719 VDD.n737 0.0405
R28684 VDD.n1720 VDD.n1719 0.0405
R28685 VDD.n1721 VDD.n1720 0.0405
R28686 VDD.n1721 VDD.n724 0.0405
R28687 VDD.n1744 VDD.n724 0.0405
R28688 VDD.n1745 VDD.n1744 0.0405
R28689 VDD.n1746 VDD.n1745 0.0405
R28690 VDD.n1746 VDD.n713 0.0405
R28691 VDD.n1772 VDD.n713 0.0405
R28692 VDD.n1773 VDD.n1772 0.0405
R28693 VDD.n1774 VDD.n701 0.0405
R28694 VDD.n1792 VDD.n701 0.0405
R28695 VDD.n1793 VDD.n1792 0.0405
R28696 VDD.n1794 VDD.n1793 0.0405
R28697 VDD.n1794 VDD.n690 0.0405
R28698 VDD.n1821 VDD.n690 0.0405
R28699 VDD.n1822 VDD.n1821 0.0405
R28700 VDD.n1823 VDD.n1822 0.0405
R28701 VDD.n1823 VDD.n681 0.0405
R28702 VDD.n1845 VDD.n681 0.0405
R28703 VDD.n1846 VDD.n1845 0.0405
R28704 VDD.n1847 VDD.n1846 0.0405
R28705 VDD.n1698 VDD.n750 0.0405
R28706 VDD.n1698 VDD.n748 0.0405
R28707 VDD.n1702 VDD.n748 0.0405
R28708 VDD.n1702 VDD.n738 0.0405
R28709 VDD.n1718 VDD.n738 0.0405
R28710 VDD.n1718 VDD.n736 0.0405
R28711 VDD.n1722 VDD.n736 0.0405
R28712 VDD.n1722 VDD.n725 0.0405
R28713 VDD.n1743 VDD.n725 0.0405
R28714 VDD.n1743 VDD.n723 0.0405
R28715 VDD.n1747 VDD.n723 0.0405
R28716 VDD.n1747 VDD.n714 0.0405
R28717 VDD.n1771 VDD.n714 0.0405
R28718 VDD.n1771 VDD.n712 0.0405
R28719 VDD.n1775 VDD.n702 0.0405
R28720 VDD.n1791 VDD.n702 0.0405
R28721 VDD.n1791 VDD.n700 0.0405
R28722 VDD.n1795 VDD.n700 0.0405
R28723 VDD.n1795 VDD.n691 0.0405
R28724 VDD.n1820 VDD.n691 0.0405
R28725 VDD.n1820 VDD.n689 0.0405
R28726 VDD.n1824 VDD.n689 0.0405
R28727 VDD.n1824 VDD.n682 0.0405
R28728 VDD.n1844 VDD.n682 0.0405
R28729 VDD.n1844 VDD.n680 0.0405
R28730 VDD.n1851 VDD.n680 0.0405
R28731 VDD.n1464 VDD.n879 0.0405
R28732 VDD.n1440 VDD.n879 0.0405
R28733 VDD.n1440 VDD.n1439 0.0405
R28734 VDD.n1439 VDD.n1438 0.0405
R28735 VDD.n1438 VDD.n917 0.0405
R28736 VDD.n1434 VDD.n917 0.0405
R28737 VDD.n1434 VDD.n1433 0.0405
R28738 VDD.n1433 VDD.n1432 0.0405
R28739 VDD.n1432 VDD.n922 0.0405
R28740 VDD.n1428 VDD.n922 0.0405
R28741 VDD.n1428 VDD.n1427 0.0405
R28742 VDD.n1427 VDD.n1426 0.0405
R28743 VDD.n1426 VDD.n927 0.0405
R28744 VDD.n1422 VDD.n927 0.0405
R28745 VDD.n1421 VDD.n1420 0.0405
R28746 VDD.n1420 VDD.n932 0.0405
R28747 VDD.n1416 VDD.n932 0.0405
R28748 VDD.n1416 VDD.n1415 0.0405
R28749 VDD.n1415 VDD.n1414 0.0405
R28750 VDD.n1414 VDD.n937 0.0405
R28751 VDD.n1410 VDD.n937 0.0405
R28752 VDD.n1410 VDD.n1409 0.0405
R28753 VDD.n1409 VDD.n1408 0.0405
R28754 VDD.n1408 VDD.n942 0.0405
R28755 VDD.n1404 VDD.n942 0.0405
R28756 VDD.n1404 VDD.n1403 0.0405
R28757 VDD.n1423 VDD.n931 0.0360676
R28758 VDD.n1774 VDD.n1773 0.0360676
R28759 VDD.n1775 VDD.n712 0.0360676
R28760 VDD.n1468 VDD.n878 0.0360676
R28761 VDD.n878 VDD.n866 0.0360676
R28762 VDD.n1490 VDD.n866 0.0360676
R28763 VDD.n1490 VDD.n864 0.0360676
R28764 VDD.n1494 VDD.n864 0.0360676
R28765 VDD.n1494 VDD.n852 0.0360676
R28766 VDD.n1514 VDD.n852 0.0360676
R28767 VDD.n1514 VDD.n849 0.0360676
R28768 VDD.n1525 VDD.n849 0.0360676
R28769 VDD.n1525 VDD.n850 0.0360676
R28770 VDD.n1521 VDD.n850 0.0360676
R28771 VDD.n1521 VDD.n1520 0.0360676
R28772 VDD.n1520 VDD.n1519 0.0360676
R28773 VDD.n1519 VDD.n823 0.0360676
R28774 VDD.n1570 VDD.n823 0.0360676
R28775 VDD.n1570 VDD.n821 0.0360676
R28776 VDD.n1574 VDD.n821 0.0360676
R28777 VDD.n1574 VDD.n810 0.0360676
R28778 VDD.n1594 VDD.n810 0.0360676
R28779 VDD.n1594 VDD.n808 0.0360676
R28780 VDD.n1598 VDD.n808 0.0360676
R28781 VDD.n1598 VDD.n797 0.0360676
R28782 VDD.n1620 VDD.n797 0.0360676
R28783 VDD.n1620 VDD.n795 0.0360676
R28784 VDD.n1624 VDD.n795 0.0360676
R28785 VDD.n1624 VDD.n784 0.0360676
R28786 VDD.n1646 VDD.n784 0.0360676
R28787 VDD.n1646 VDD.n781 0.0360676
R28788 VDD.n1651 VDD.n781 0.0360676
R28789 VDD.n1651 VDD.n782 0.0360676
R28790 VDD.n782 VDD.n768 0.0360676
R28791 VDD.n1680 VDD.n768 0.0360676
R28792 VDD.n1680 VDD.n766 0.0360676
R28793 VDD.n1467 VDD.n1466 0.0360676
R28794 VDD.n1466 VDD.n865 0.0360676
R28795 VDD.n1491 VDD.n865 0.0360676
R28796 VDD.n1492 VDD.n1491 0.0360676
R28797 VDD.n1493 VDD.n1492 0.0360676
R28798 VDD.n1493 VDD.n851 0.0360676
R28799 VDD.n1515 VDD.n851 0.0360676
R28800 VDD.n1516 VDD.n1515 0.0360676
R28801 VDD.n1524 VDD.n1516 0.0360676
R28802 VDD.n1524 VDD.n1523 0.0360676
R28803 VDD.n1523 VDD.n1522 0.0360676
R28804 VDD.n1522 VDD.n1517 0.0360676
R28805 VDD.n1518 VDD.n1517 0.0360676
R28806 VDD.n1518 VDD.n822 0.0360676
R28807 VDD.n1571 VDD.n822 0.0360676
R28808 VDD.n1572 VDD.n1571 0.0360676
R28809 VDD.n1573 VDD.n1572 0.0360676
R28810 VDD.n1573 VDD.n809 0.0360676
R28811 VDD.n1595 VDD.n809 0.0360676
R28812 VDD.n1596 VDD.n1595 0.0360676
R28813 VDD.n1597 VDD.n1596 0.0360676
R28814 VDD.n1597 VDD.n796 0.0360676
R28815 VDD.n1621 VDD.n796 0.0360676
R28816 VDD.n1622 VDD.n1621 0.0360676
R28817 VDD.n1623 VDD.n1622 0.0360676
R28818 VDD.n1623 VDD.n783 0.0360676
R28819 VDD.n1647 VDD.n783 0.0360676
R28820 VDD.n1648 VDD.n1647 0.0360676
R28821 VDD.n1650 VDD.n1648 0.0360676
R28822 VDD.n1650 VDD.n1649 0.0360676
R28823 VDD.n1649 VDD.n767 0.0360676
R28824 VDD.n1681 VDD.n767 0.0360676
R28825 VDD.n1682 VDD.n1681 0.0360676
R28826 VDD.n1422 VDD.n1421 0.0360676
R28827 VDD.n1308 VDD.n947 0.0360676
R28828 VDD.n1309 VDD.n1308 0.0360676
R28829 VDD.n1310 VDD.n1309 0.0360676
R28830 VDD.n1311 VDD.n1310 0.0360676
R28831 VDD.n1325 VDD.n1311 0.0360676
R28832 VDD.n1326 VDD.n1325 0.0360676
R28833 VDD.n1327 VDD.n1326 0.0360676
R28834 VDD.n1343 VDD.n1327 0.0360676
R28835 VDD.n1344 VDD.n1343 0.0360676
R28836 VDD.n1356 VDD.n1344 0.0360676
R28837 VDD.n1356 VDD.n1355 0.0360676
R28838 VDD.n1355 VDD.n1352 0.0360676
R28839 VDD.n1352 VDD.n1351 0.0360676
R28840 VDD.n1351 VDD.n1348 0.0360676
R28841 VDD.n1348 VDD.n1347 0.0360676
R28842 VDD.n1347 VDD.n1345 0.0360676
R28843 VDD.n1345 VDD.n600 0.0360676
R28844 VDD.n601 VDD.n600 0.0360676
R28845 VDD.n618 VDD.n601 0.0360676
R28846 VDD.n619 VDD.n618 0.0360676
R28847 VDD.n620 VDD.n619 0.0360676
R28848 VDD.n621 VDD.n620 0.0360676
R28849 VDD.n638 VDD.n621 0.0360676
R28850 VDD.n639 VDD.n638 0.0360676
R28851 VDD.n640 VDD.n639 0.0360676
R28852 VDD.n641 VDD.n640 0.0360676
R28853 VDD.n659 VDD.n641 0.0360676
R28854 VDD.n660 VDD.n659 0.0360676
R28855 VDD.n663 VDD.n660 0.0360676
R28856 VDD.n664 VDD.n663 0.0360676
R28857 VDD.n665 VDD.n664 0.0360676
R28858 VDD.n666 VDD.n665 0.0360676
R28859 VDD.n1848 VDD.n666 0.0360676
R28860 VDD.n1307 VDD.n948 0.0360676
R28861 VDD.n1307 VDD.n1306 0.0360676
R28862 VDD.n1383 VDD.n1306 0.0360676
R28863 VDD.n1383 VDD.n1382 0.0360676
R28864 VDD.n1382 VDD.n1312 0.0360676
R28865 VDD.n1371 VDD.n1312 0.0360676
R28866 VDD.n1371 VDD.n1370 0.0360676
R28867 VDD.n1370 VDD.n1328 0.0360676
R28868 VDD.n1358 VDD.n1328 0.0360676
R28869 VDD.n1358 VDD.n1357 0.0360676
R28870 VDD.n1354 VDD.n1353 0.0360676
R28871 VDD.n1350 VDD.n1349 0.0360676
R28872 VDD.n1346 VDD.n599 0.0360676
R28873 VDD.n1923 VDD.n599 0.0360676
R28874 VDD.n1923 VDD.n1922 0.0360676
R28875 VDD.n1922 VDD.n602 0.0360676
R28876 VDD.n617 VDD.n602 0.0360676
R28877 VDD.n1911 VDD.n617 0.0360676
R28878 VDD.n1911 VDD.n1910 0.0360676
R28879 VDD.n1910 VDD.n622 0.0360676
R28880 VDD.n637 VDD.n622 0.0360676
R28881 VDD.n1898 VDD.n637 0.0360676
R28882 VDD.n1898 VDD.n1897 0.0360676
R28883 VDD.n1897 VDD.n642 0.0360676
R28884 VDD.n661 VDD.n642 0.0360676
R28885 VDD.n662 VDD.n661 0.0360676
R28886 VDD.n662 VDD.n658 0.0360676
R28887 VDD.n1876 VDD.n658 0.0360676
R28888 VDD.n1876 VDD.n1875 0.0360676
R28889 VDD.n1875 VDD.n667 0.0360676
R28890 VDD VDD.n296 0.0358992
R28891 VDD VDD.n291 0.0358992
R28892 VDD.n2044 VDD 0.0358992
R28893 VDD.n2035 VDD 0.0358992
R28894 VDD.n285 VDD 0.0355649
R28895 VDD.n2025 VDD 0.0355649
R28896 VDD.n582 VDD.n577 0.0262169
R28897 VDD.n1463 VDD.n877 0.0234189
R28898 VDD.n1683 VDD.n749 0.0234189
R28899 VDD.n1684 VDD.n750 0.0234189
R28900 VDD.n1465 VDD.n1464 0.0234189
R28901 VDD.n75 VDD.n74 0.023342
R28902 VDD.n1401 VDD.n946 0.0233108
R28903 VDD.n1849 VDD.n1847 0.0233108
R28904 VDD.n1851 VDD.n1850 0.0233108
R28905 VDD.n1403 VDD.n1402 0.0233108
R28906 VDD.n1468 VDD.n877 0.0227703
R28907 VDD.n1467 VDD.n1465 0.0227703
R28908 VDD.n1402 VDD.n947 0.0227703
R28909 VDD.n1401 VDD.n948 0.0227703
R28910 VDD.n2046 VDD 0.0221393
R28911 VDD.n2034 VDD 0.0221393
R28912 VDD VDD.n2050 0.0221393
R28913 VDD.n74 VDD.n73 0.0219014
R28914 VDD.n1443 VDD.n911 0.0188784
R28915 VDD.n1045 VDD.n915 0.0188784
R28916 VDD.n1054 VDD.n1053 0.0188784
R28917 VDD.n1063 VDD.n1062 0.0188784
R28918 VDD.n1070 VDD.n1069 0.0188784
R28919 VDD.n1096 VDD.n1095 0.0188784
R28920 VDD.n1104 VDD.n1103 0.0188784
R28921 VDD.n1111 VDD.n1110 0.0188784
R28922 VDD.n1126 VDD.n1012 0.0188784
R28923 VDD.n1129 VDD.n1128 0.0188784
R28924 VDD.n1143 VDD.n1005 0.0188784
R28925 VDD.n1153 VDD.n1152 0.0188784
R28926 VDD.n1162 VDD.n1161 0.0188784
R28927 VDD.n1171 VDD.n1170 0.0188784
R28928 VDD.n1180 VDD.n1179 0.0188784
R28929 VDD.n1187 VDD.n1186 0.0188784
R28930 VDD.n1198 VDD.n1196 0.0188784
R28931 VDD.n1212 VDD.n981 0.0188784
R28932 VDD.n1228 VDD.n1227 0.0188784
R28933 VDD.n1243 VDD.n969 0.0188784
R28934 VDD.n1246 VDD.n1245 0.0188784
R28935 VDD.n1254 VDD.n1253 0.0188784
R28936 VDD.n1268 VDD.n961 0.0188784
R28937 VDD.n1400 VDD.n950 0.0188784
R28938 VDD.n1300 VDD.n1299 0.0188784
R28939 VDD.n1390 VDD.n1389 0.0188784
R28940 VDD.n1386 VDD.n1385 0.0188784
R28941 VDD.n759 VDD.n752 0.0188784
R28942 VDD.n757 VDD.n747 0.0188784
R28943 VDD.n1707 VDD.n1704 0.0188784
R28944 VDD.n1705 VDD.n739 0.0188784
R28945 VDD.n1716 VDD.n741 0.0188784
R28946 VDD.n1730 VDD.n1729 0.0188784
R28947 VDD.n1732 VDD.n726 0.0188784
R28948 VDD.n1741 VDD.n728 0.0188784
R28949 VDD.n1749 VDD.n722 0.0188784
R28950 VDD.n1754 VDD.n720 0.0188784
R28951 VDD.n1757 VDD.n1756 0.0188784
R28952 VDD.n1769 VDD.n716 0.0188784
R28953 VDD.n1765 VDD.n711 0.0188784
R28954 VDD.n1780 VDD.n1777 0.0188784
R28955 VDD.n1778 VDD.n703 0.0188784
R28956 VDD.n1789 VDD.n705 0.0188784
R28957 VDD.n1797 VDD.n699 0.0188784
R28958 VDD.n1802 VDD.n697 0.0188784
R28959 VDD.n1818 VDD.n693 0.0188784
R28960 VDD.n1813 VDD.n688 0.0188784
R28961 VDD.n1829 VDD.n1826 0.0188784
R28962 VDD.n1827 VDD.n683 0.0188784
R28963 VDD.n1842 VDD.n684 0.0188784
R28964 VDD.n1925 VDD.n596 0.0188784
R28965 VDD.n603 VDD.n598 0.0188784
R28966 VDD.n1920 VDD.n604 0.0188784
R28967 VDD.n614 VDD.n613 0.0188784
R28968 VDD.n886 VDD.n876 0.0188784
R28969 VDD.n1471 VDD.n1470 0.0188784
R28970 VDD.n1480 VDD.n1479 0.0188784
R28971 VDD.n1482 VDD.n867 0.0188784
R28972 VDD.n1563 VDD.n820 0.0188784
R28973 VDD.n1579 VDD.n1576 0.0188784
R28974 VDD.n1577 VDD.n811 0.0188784
R28975 VDD.n1592 VDD.n813 0.0188784
R28976 VDD.n1461 VDD.n882 0.0187703
R28977 VDD.n911 VDD.n910 0.0187703
R28978 VDD.n1081 VDD.n1079 0.0187703
R28979 VDD.n1095 VDD.n1024 0.0187703
R28980 VDD.n1144 VDD.n1143 0.0187703
R28981 VDD.n1213 VDD.n1212 0.0187703
R28982 VDD.n1221 VDD.n1220 0.0187703
R28983 VDD.n1269 VDD.n1268 0.0187703
R28984 VDD.n1278 VDD.n1277 0.0187703
R28985 VDD.n1380 VDD.n1313 0.0187703
R28986 VDD.n1373 VDD.n1323 0.0187703
R28987 VDD.n1329 VDD.n1324 0.0187703
R28988 VDD.n1368 VDD.n1330 0.0187703
R28989 VDD.n1342 VDD.n1341 0.0187703
R28990 VDD.n1360 VDD.n583 0.0187703
R28991 VDD.n1688 VDD.n751 0.0187703
R28992 VDD.n1696 VDD.n752 0.0187703
R28993 VDD.n1724 VDD.n735 0.0187703
R28994 VDD.n1729 VDD.n733 0.0187703
R28995 VDD.n1757 VDD.n715 0.0187703
R28996 VDD.n1803 VDD.n1802 0.0187703
R28997 VDD.n1805 VDD.n692 0.0187703
R28998 VDD.n1837 VDD.n684 0.0187703
R28999 VDD.n1853 VDD.n678 0.0187703
R29000 VDD.n623 VDD.n616 0.0187703
R29001 VDD.n1908 VDD.n624 0.0187703
R29002 VDD.n634 VDD.n633 0.0187703
R29003 VDD.n1901 VDD.n1900 0.0187703
R29004 VDD.n643 VDD.n636 0.0187703
R29005 VDD.n1895 VDD.n644 0.0187703
R29006 VDD.n1891 VDD.n1890 0.0187703
R29007 VDD.n1887 VDD.n1886 0.0187703
R29008 VDD.n1883 VDD.n1882 0.0187703
R29009 VDD.n1879 VDD.n1878 0.0187703
R29010 VDD.n668 VDD.n657 0.0187703
R29011 VDD.n1873 VDD.n669 0.0187703
R29012 VDD.n1496 VDD.n863 0.0187703
R29013 VDD.n1504 VDD.n856 0.0187703
R29014 VDD.n1506 VDD.n853 0.0187703
R29015 VDD.n1512 VDD.n854 0.0187703
R29016 VDD.n1528 VDD.n1527 0.0187703
R29017 VDD.n848 VDD.n846 0.0187703
R29018 VDD.n1538 VDD.n1537 0.0187703
R29019 VDD.n1542 VDD.n1541 0.0187703
R29020 VDD.n1546 VDD.n1545 0.0187703
R29021 VDD.n1551 VDD.n1550 0.0187703
R29022 VDD.n1553 VDD.n824 0.0187703
R29023 VDD.n1568 VDD.n825 0.0187703
R29024 VDD.n1604 VDD.n1600 0.0187703
R29025 VDD.n1602 VDD.n798 0.0187703
R29026 VDD.n1618 VDD.n799 0.0187703
R29027 VDD.n1612 VDD.n794 0.0187703
R29028 VDD.n1630 VDD.n1629 0.0187703
R29029 VDD.n1627 VDD.n785 0.0187703
R29030 VDD.n1644 VDD.n786 0.0187703
R29031 VDD.n1639 VDD.n780 0.0187703
R29032 VDD.n1654 VDD.n1653 0.0187703
R29033 VDD.n1667 VDD.n1664 0.0187703
R29034 VDD.n1665 VDD.n769 0.0187703
R29035 VDD.n1678 VDD.n770 0.0187703
R29036 VDD.n1357 VDD.n590 0.0186443
R29037 VDD.n1353 VDD.n589 0.0186443
R29038 VDD.n1349 VDD.n588 0.0186443
R29039 VDD.n1354 VDD.n590 0.0186443
R29040 VDD.n1350 VDD.n589 0.0186443
R29041 VDD.n1346 VDD.n588 0.0186443
R29042 VDD.n1442 VDD.n915 0.0185541
R29043 VDD.n1253 VDD.n944 0.0185541
R29044 VDD.n758 VDD.n757 0.0185541
R29045 VDD.n1843 VDD.n683 0.0185541
R29046 VDD.n1381 VDD.n1305 0.0184459
R29047 VDD.n1913 VDD.n1912 0.0184459
R29048 VDD.n1488 VDD.n868 0.0184459
R29049 VDD.n1599 VDD.n807 0.0184459
R29050 VDD.n1152 VDD.n929 0.0182297
R29051 VDD.n1770 VDD.n1769 0.0182297
R29052 VDD.n1384 VDD.n1305 0.0181216
R29053 VDD.n1913 VDD.n615 0.0181216
R29054 VDD.n1489 VDD.n1488 0.0181216
R29055 VDD.n812 VDD.n807 0.0181216
R29056 VDD.n1081 VDD.n1080 0.0175811
R29057 VDD.n1220 VDD.n938 0.0175811
R29058 VDD.n1724 VDD.n1723 0.0175811
R29059 VDD.n1805 VDD.n1804 0.0175811
R29060 VDD.n1322 VDD.n1313 0.0173649
R29061 VDD.n1909 VDD.n623 0.0173649
R29062 VDD.n1496 VDD.n1495 0.0173649
R29063 VDD.n1604 VDD.n1603 0.0173649
R29064 VDD.n1386 VDD.n1303 0.0170405
R29065 VDD.n613 VDD.n611 0.0170405
R29066 VDD.n1482 VDD.n1481 0.0170405
R29067 VDD.n1593 VDD.n1592 0.0170405
R29068 VDD.n1103 VDD.n923 0.0167162
R29069 VDD.n1198 VDD.n1197 0.0167162
R29070 VDD.n1732 VDD.n1731 0.0167162
R29071 VDD.n1797 VDD.n1796 0.0167162
R29072 VDD.n1373 VDD.n1372 0.0162838
R29073 VDD.n631 VDD.n624 0.0162838
R29074 VDD.n1505 VDD.n1504 0.0162838
R29075 VDD.n1619 VDD.n798 0.0162838
R29076 VDD.n1128 VDD.n928 0.0159595
R29077 VDD.n1170 VDD.n994 0.0159595
R29078 VDD.n1390 VDD.n1302 0.0159595
R29079 VDD.n1755 VDD.n1754 0.0159595
R29080 VDD.n1777 VDD.n1776 0.0159595
R29081 VDD.n1921 VDD.n1920 0.0159595
R29082 VDD.n1479 VDD.n870 0.0159595
R29083 VDD.n1578 VDD.n1577 0.0159595
R29084 VDD.n909 VDD.n882 0.0157432
R29085 VDD.n1278 VDD.n945 0.0157432
R29086 VDD.n1697 VDD.n751 0.0157432
R29087 VDD.n1836 VDD.n678 0.0157432
R29088 VDD.n1053 VDD.n1037 0.0152027
R29089 VDD.n1245 VDD.n943 0.0152027
R29090 VDD.n1369 VDD.n1329 0.0152027
R29091 VDD.n1704 VDD.n1703 0.0152027
R29092 VDD.n1829 VDD.n1828 0.0152027
R29093 VDD.n635 VDD.n634 0.0152027
R29094 VDD.n1513 VDD.n853 0.0152027
R29095 VDD.n1611 VDD.n799 0.0152027
R29096 VDD.n1161 VDD.n930 0.0148784
R29097 VDD.n1299 VDD.n1298 0.0148784
R29098 VDD.n1765 VDD.n1764 0.0148784
R29099 VDD.n1924 VDD.n598 0.0148784
R29100 VDD.n1470 VDD.n1469 0.0148784
R29101 VDD.n1576 VDD.n1575 0.0148784
R29102 VDD.n455 VDD.n423 0.0148556
R29103 VDD.n511 VDD.n510 0.0148556
R29104 VDD.n1069 VDD.n920 0.0141216
R29105 VDD.n1227 VDD.n939 0.0141216
R29106 VDD.n1340 VDD.n1330 0.0141216
R29107 VDD.n741 VDD.n740 0.0141216
R29108 VDD.n1819 VDD.n1818 0.0141216
R29109 VDD.n1900 VDD.n1899 0.0141216
R29110 VDD.n854 VDD.n845 0.0141216
R29111 VDD.n1625 VDD.n794 0.0141216
R29112 VDD.n596 VDD.n584 0.0137973
R29113 VDD.n673 VDD.n672 0.0137973
R29114 VDD.n1563 VDD.n1562 0.0137973
R29115 VDD.n1685 VDD.n763 0.0137973
R29116 VDD.n1684 VDD.n766 0.0137973
R29117 VDD.n1683 VDD.n1682 0.0137973
R29118 VDD.n1849 VDD.n1848 0.0137973
R29119 VDD.n1850 VDD.n667 0.0137973
R29120 VDD.n1869 VDD.n1868 0.0134381
R29121 VDD.n1110 VDD.n924 0.0133649
R29122 VDD.n1186 VDD.n935 0.0133649
R29123 VDD.n1742 VDD.n1741 0.0133649
R29124 VDD.n705 VDD.n704 0.0133649
R29125 VDD.n1359 VDD.n1342 0.0130405
R29126 VDD.n1896 VDD.n643 0.0130405
R29127 VDD.n1527 VDD.n1526 0.0130405
R29128 VDD.n1629 VDD.n1628 0.0130405
R29129 VDD.n1874 VDD.n1873 0.0128243
R29130 VDD.n1569 VDD.n1568 0.0128243
R29131 VDD.n1679 VDD.n1678 0.0128243
R29132 VDD.n2047 VDD.n2046 0.0126721
R29133 VDD.n2034 VDD.n2021 0.0126721
R29134 VDD.n2050 VDD.n2049 0.0126721
R29135 VDD.n1127 VDD.n1126 0.0126081
R29136 VDD.n1179 VDD.n933 0.0126081
R29137 VDD.n1749 VDD.n1748 0.0126081
R29138 VDD.n1779 VDD.n1778 0.0126081
R29139 VDD.n1462 VDD.n881 0.0123919
R29140 VDD.n1276 VDD.n949 0.0123919
R29141 VDD.n1687 VDD.n1686 0.0123919
R29142 VDD.n1852 VDD.n679 0.0123919
R29143 VDD.n650 VDD.n644 0.0119595
R29144 VDD.n846 VDD.n838 0.0119595
R29145 VDD.n1645 VDD.n785 0.0119595
R29146 VDD.n1062 VDD.n918 0.0118514
R29147 VDD.n1244 VDD.n1243 0.0118514
R29148 VDD.n1706 VDD.n1705 0.0118514
R29149 VDD.n1825 VDD.n688 0.0118514
R29150 VDD.n1877 VDD.n657 0.0117432
R29151 VDD.n1553 VDD.n1552 0.0117432
R29152 VDD.n1666 VDD.n1665 0.0117432
R29153 VDD.n1673 VDD.n761 0.0116588
R29154 VDD.n886 VDD.n881 0.011527
R29155 VDD.n1686 VDD.n1685 0.011527
R29156 VDD.n1400 VDD.n949 0.0114189
R29157 VDD.n679 VDD.n673 0.0114189
R29158 VDD.n1476 VDD.n860 0.0109762
R29159 VDD.n1501 VDD.n1500 0.0109762
R29160 VDD.n1531 VDD.n842 0.0109762
R29161 VDD.n1534 VDD.n1532 0.0109762
R29162 VDD.n1533 VDD.n829 0.0109762
R29163 VDD.n1558 VDD.n1557 0.0109762
R29164 VDD.n1583 VDD.n817 0.0109762
R29165 VDD.n1584 VDD.n804 0.0109762
R29166 VDD.n1609 VDD.n1608 0.0109762
R29167 VDD.n1633 VDD.n791 0.0109762
R29168 VDD.n1635 VDD.n1634 0.0109762
R29169 VDD.n1692 VDD.n1691 0.0109762
R29170 VDD.n1692 VDD.n743 0.0109762
R29171 VDD.n1710 VDD.n743 0.0109762
R29172 VDD.n1711 VDD.n1710 0.0109762
R29173 VDD.n1712 VDD.n1711 0.0109762
R29174 VDD.n1712 VDD.n730 0.0109762
R29175 VDD.n1735 VDD.n730 0.0109762
R29176 VDD.n1736 VDD.n1735 0.0109762
R29177 VDD.n1737 VDD.n1736 0.0109762
R29178 VDD.n1737 VDD.n718 0.0109762
R29179 VDD.n1760 VDD.n718 0.0109762
R29180 VDD.n1761 VDD.n707 0.0109762
R29181 VDD.n1783 VDD.n707 0.0109762
R29182 VDD.n1784 VDD.n1783 0.0109762
R29183 VDD.n1785 VDD.n1784 0.0109762
R29184 VDD.n1785 VDD.n695 0.0109762
R29185 VDD.n1808 VDD.n695 0.0109762
R29186 VDD.n1809 VDD.n1808 0.0109762
R29187 VDD.n1809 VDD.n686 0.0109762
R29188 VDD.n1832 VDD.n686 0.0109762
R29189 VDD.n1833 VDD.n1832 0.0109762
R29190 VDD.n1833 VDD.n676 0.0109762
R29191 VDD.n1856 VDD.n676 0.0109762
R29192 VDD.n1318 VDD.n1316 0.0109762
R29193 VDD.n1377 VDD.n1376 0.0109762
R29194 VDD.n1364 VDD.n1319 0.0109762
R29195 VDD.n1363 VDD.n1337 0.0109762
R29196 VDD.n1335 VDD.n594 0.0109762
R29197 VDD.n1931 VDD.n1930 0.0109762
R29198 VDD.n1928 VDD.n595 0.0109762
R29199 VDD.n1917 VDD.n1916 0.0109762
R29200 VDD.n1905 VDD.n608 0.0109762
R29201 VDD.n1904 VDD.n628 0.0109762
R29202 VDD.n1861 VDD.n1860 0.0109762
R29203 VDD.n1863 VDD.n1862 0.0109762
R29204 VDD.n1868 VDD.n1867 0.0109762
R29205 VDD.n1476 VDD.n1475 0.01095
R29206 VDD.n1500 VDD.n860 0.01095
R29207 VDD.n1501 VDD.n842 0.01095
R29208 VDD.n1532 VDD.n1531 0.01095
R29209 VDD.n1534 VDD.n1533 0.01095
R29210 VDD.n1557 VDD.n829 0.01095
R29211 VDD.n1558 VDD.n817 0.01095
R29212 VDD.n1584 VDD.n1583 0.01095
R29213 VDD.n1608 VDD.n804 0.01095
R29214 VDD.n1609 VDD.n791 0.01095
R29215 VDD.n1634 VDD.n1633 0.01095
R29216 VDD.n1636 VDD.n1635 0.01095
R29217 VDD.n1761 VDD.n1760 0.01095
R29218 VDD.n1857 VDD.n1856 0.01095
R29219 VDD.n1377 VDD.n1318 0.01095
R29220 VDD.n1376 VDD.n1319 0.01095
R29221 VDD.n1364 VDD.n1363 0.01095
R29222 VDD.n1337 VDD.n1335 0.01095
R29223 VDD.n1931 VDD.n594 0.01095
R29224 VDD.n1930 VDD.n1928 0.01095
R29225 VDD.n1917 VDD.n595 0.01095
R29226 VDD.n1916 VDD.n608 0.01095
R29227 VDD.n1905 VDD.n1904 0.01095
R29228 VDD.n1860 VDD.n628 0.01095
R29229 VDD.n1862 VDD.n1861 0.01095
R29230 VDD.n1867 VDD.n1863 0.01095
R29231 VDD.n1890 VDD.n651 0.0108784
R29232 VDD.n1538 VDD.n836 0.0108784
R29233 VDD.n1638 VDD.n786 0.0108784
R29234 VDD.n1063 VDD.n919 0.0107703
R29235 VDD.n969 VDD.n940 0.0107703
R29236 VDD.n1717 VDD.n739 0.0107703
R29237 VDD.n1813 VDD.n1812 0.0107703
R29238 VDD.n1879 VDD.n655 0.0106622
R29239 VDD.n1550 VDD.n832 0.0106622
R29240 VDD.n1664 VDD.n776 0.0106622
R29241 VDD.n1691 VDD.n761 0.0106095
R29242 VDD.n1012 VDD.n925 0.0100135
R29243 VDD.n1180 VDD.n934 0.0100135
R29244 VDD.n727 VDD.n722 0.0100135
R29245 VDD.n1790 VDD.n703 0.0100135
R29246 VDD.n1886 VDD.n653 0.0097973
R29247 VDD.n1542 VDD.n834 0.0097973
R29248 VDD.n1652 VDD.n780 0.0097973
R29249 VDD.n1674 VDD.n1673 0.00967266
R29250 VDD.n1883 VDD.n653 0.00958108
R29251 VDD.n1545 VDD.n834 0.00958108
R29252 VDD.n1654 VDD.n1652 0.00958108
R29253 VDD.n1111 VDD.n925 0.00925676
R29254 VDD.n1187 VDD.n934 0.00925676
R29255 VDD.n728 VDD.n727 0.00925676
R29256 VDD.n1790 VDD.n1789 0.00925676
R29257 VDD.n1557 VDD.n828 0.00880612
R29258 VDD.n1882 VDD.n655 0.00871622
R29259 VDD.n1546 VDD.n832 0.00871622
R29260 VDD.n1653 VDD.n776 0.00871622
R29261 VDD.n562 VDD 0.00859195
R29262 VDD.n580 VDD.n577 0.00853653
R29263 VDD.n580 VDD.n579 0.00853653
R29264 VDD.n1070 VDD.n919 0.0085
R29265 VDD.n1228 VDD.n940 0.0085
R29266 VDD.n1717 VDD.n1716 0.0085
R29267 VDD.n1812 VDD.n693 0.0085
R29268 VDD.n1887 VDD.n651 0.0085
R29269 VDD.n1541 VDD.n836 0.0085
R29270 VDD.n1639 VDD.n1638 0.0085
R29271 VDD.n1316 VDD.n1297 0.00809524
R29272 VDD.n1672 VDD.n1671 0.00778095
R29273 VDD.n1934 VDD.n583 0.00763514
R29274 VDD.n1878 VDD.n1877 0.00763514
R29275 VDD.n1552 VDD.n1551 0.00763514
R29276 VDD.n1667 VDD.n1666 0.00763514
R29277 VDD.n1054 VDD.n918 0.00741892
R29278 VDD.n1246 VDD.n1244 0.00741892
R29279 VDD.n1707 VDD.n1706 0.00741892
R29280 VDD.n1826 VDD.n1825 0.00741892
R29281 VDD.n1891 VDD.n650 0.00741892
R29282 VDD.n1537 VDD.n838 0.00741892
R29283 VDD.n1645 VDD.n1644 0.00741892
R29284 VDD.n1636 VDD.n778 0.00725714
R29285 VDD.n1674 VDD.n1672 0.00707381
R29286 VDD.n1462 VDD.n1461 0.00698649
R29287 VDD.n1277 VDD.n1276 0.00698649
R29288 VDD.n1688 VDD.n1687 0.00698649
R29289 VDD.n1853 VDD.n1852 0.00698649
R29290 VDD.n1475 VDD.n874 0.00696162
R29291 VDD.n1857 VDD.n675 0.00691667
R29292 VDD.n1129 VDD.n1127 0.00666216
R29293 VDD.n1171 VDD.n933 0.00666216
R29294 VDD.n1748 VDD.n720 0.00666216
R29295 VDD.n1780 VDD.n1779 0.00666216
R29296 VDD.n1927 VDD.n585 0.00660407
R29297 VDD.n1874 VDD.n668 0.00655405
R29298 VDD.n1569 VDD.n824 0.00655405
R29299 VDD.n1679 VDD.n769 0.00655405
R29300 VDD.n593 VDD.n592 0.00634975
R29301 VDD.n1360 VDD.n1359 0.00633784
R29302 VDD.n1896 VDD.n1895 0.00633784
R29303 VDD.n1526 VDD.n848 0.00633784
R29304 VDD.n1628 VDD.n1627 0.00633784
R29305 VDD.n1933 VDD.n1932 0.00613116
R29306 VDD.n1104 VDD.n924 0.00590541
R29307 VDD.n1196 VDD.n935 0.00590541
R29308 VDD.n1742 VDD.n726 0.00590541
R29309 VDD.n704 VDD.n699 0.00590541
R29310 VDD.n1583 VDD.n816 0.00588776
R29311 VDD.n1475 VDD.n873 0.00588776
R29312 VDD.n1336 VDD.n591 0.00581903
R29313 VDD.n1933 VDD.n593 0.00567741
R29314 VDD.n1932 VDD.n586 0.00556475
R29315 VDD.n672 VDD.n669 0.00547297
R29316 VDD.n1562 VDD.n825 0.00547297
R29317 VDD.n770 VDD.n763 0.00547297
R29318 VDD.n1929 VDD.n586 0.00527728
R29319 VDD.n1341 VDD.n1340 0.00525676
R29320 VDD.n1899 VDD.n636 0.00525676
R29321 VDD.n1528 VDD.n845 0.00525676
R29322 VDD.n1630 VDD.n1625 0.00525676
R29323 VDD.n1079 VDD.n920 0.00514865
R29324 VDD.n1221 VDD.n939 0.00514865
R29325 VDD.n740 VDD.n735 0.00514865
R29326 VDD.n1819 VDD.n692 0.00514865
R29327 VDD.n1334 VDD.n591 0.00500085
R29328 VDD.n1934 VDD.n584 0.00460811
R29329 VDD.n1334 VDD.n592 0.00449225
R29330 VDD.n1869 VDD.n1859 0.00440238
R29331 VDD.n1153 VDD.n930 0.00439189
R29332 VDD.n1298 VDD.n950 0.00439189
R29333 VDD.n1764 VDD.n716 0.00439189
R29334 VDD.n1925 VDD.n1924 0.00439189
R29335 VDD.n1469 VDD.n876 0.00439189
R29336 VDD.n1575 VDD.n820 0.00439189
R29337 VDD.n1689 VDD.n762 0.00425921
R29338 VDD.n1695 VDD.n753 0.00425921
R29339 VDD.n746 VDD.n745 0.00425921
R29340 VDD.n1715 VDD.n1714 0.00425921
R29341 VDD.n1728 VDD.n731 0.00425921
R29342 VDD.n1733 VDD.n732 0.00425921
R29343 VDD.n1740 VDD.n1739 0.00425921
R29344 VDD.n1750 VDD.n721 0.00425921
R29345 VDD.n1768 VDD.n1767 0.00425921
R29346 VDD.n710 VDD.n709 0.00425921
R29347 VDD.n1788 VDD.n1787 0.00425921
R29348 VDD.n1798 VDD.n698 0.00425921
R29349 VDD.n1801 VDD.n1800 0.00425921
R29350 VDD.n1817 VDD.n1816 0.00425921
R29351 VDD.n1814 VDD.n1811 0.00425921
R29352 VDD.n1838 VDD.n677 0.00425921
R29353 VDD.n1854 VDD.n671 0.00425921
R29354 VDD.n1387 VDD.n1304 0.00425921
R29355 VDD.n1379 VDD.n1314 0.00425921
R29356 VDD.n1320 VDD.n1315 0.00425921
R29357 VDD.n1374 VDD.n1321 0.00425921
R29358 VDD.n1339 VDD.n587 0.00425921
R29359 VDD.n1927 VDD.n1926 0.00425921
R29360 VDD.n612 VDD.n609 0.00425921
R29361 VDD.n1914 VDD.n610 0.00425921
R29362 VDD.n1907 VDD.n626 0.00425921
R29363 VDD.n632 VDD.n627 0.00425921
R29364 VDD.n1893 VDD.n1892 0.00425921
R29365 VDD.n1889 VDD.n1888 0.00425921
R29366 VDD.n1885 VDD.n1884 0.00425921
R29367 VDD.n1881 VDD.n1880 0.00425921
R29368 VDD.n1540 VDD.n1539 0.00425921
R29369 VDD.n1544 VDD.n1543 0.00425921
R29370 VDD.n1641 VDD.n1640 0.00425921
R29371 VDD.n1655 VDD.n779 0.00425921
R29372 VDD.n1661 VDD.n1659 0.00424524
R29373 VDD.n1695 VDD.n1694 0.0042371
R29374 VDD.n760 VDD.n756 0.0042371
R29375 VDD.n754 VDD.n744 0.0042371
R29376 VDD.n1708 VDD.n746 0.0042371
R29377 VDD.n1725 VDD.n734 0.0042371
R29378 VDD.n1728 VDD.n1727 0.0042371
R29379 VDD.n1751 VDD.n1750 0.0042371
R29380 VDD.n1753 VDD.n719 0.0042371
R29381 VDD.n1758 VDD.n717 0.0042371
R29382 VDD.n1768 VDD.n717 0.0042371
R29383 VDD.n1767 VDD.n1766 0.0042371
R29384 VDD.n1762 VDD.n708 0.0042371
R29385 VDD.n1781 VDD.n710 0.0042371
R29386 VDD.n1801 VDD.n696 0.0042371
R29387 VDD.n1806 VDD.n694 0.0042371
R29388 VDD.n1811 VDD.n687 0.0042371
R29389 VDD.n1830 VDD.n685 0.0042371
R29390 VDD.n1841 VDD.n1835 0.0042371
R29391 VDD.n1839 VDD.n1838 0.0042371
R29392 VDD.n1392 VDD.n1391 0.0042371
R29393 VDD.n1388 VDD.n1387 0.0042371
R29394 VDD.n1331 VDD.n1321 0.0042371
R29395 VDD.n1367 VDD.n1366 0.0042371
R29396 VDD.n1338 VDD.n1333 0.0042371
R29397 VDD.n1361 VDD.n1339 0.0042371
R29398 VDD.n1926 VDD.n597 0.0042371
R29399 VDD.n1919 VDD.n606 0.0042371
R29400 VDD.n612 VDD.n607 0.0042371
R29401 VDD.n632 VDD.n629 0.0042371
R29402 VDD.n1902 VDD.n630 0.0042371
R29403 VDD.n647 VDD.n646 0.0042371
R29404 VDD.n1894 VDD.n1893 0.0042371
R29405 VDD.n1880 VDD.n656 0.0042371
R29406 VDD.n1865 VDD.n1864 0.0042371
R29407 VDD.n1872 VDD.n1871 0.0042371
R29408 VDD.n1871 VDD.n1870 0.0042371
R29409 VDD.n1483 VDD.n869 0.0042371
R29410 VDD.n1511 VDD.n843 0.0042371
R29411 VDD.n1529 VDD.n844 0.0042371
R29412 VDD.n1567 VDD.n1566 0.0042371
R29413 VDD.n1591 VDD.n1586 0.0042371
R29414 VDD.n1613 VDD.n792 0.0042371
R29415 VDD.n1631 VDD.n793 0.0042371
R29416 VDD.n773 VDD.n772 0.0042371
R29417 VDD.n1677 VDD.n1676 0.0042371
R29418 VDD.n1398 VDD.n1397 0.00423273
R29419 VDD.n1566 VDD.n1565 0.00423268
R29420 VDD.n1293 VDD.n1292 0.00422178
R29421 VDD.n896 VDD.n895 0.00422178
R29422 VDD.n1658 VDD.n778 0.00421905
R29423 VDD.n1929 VDD.n585 0.00421586
R29424 VDD.n1369 VDD.n1368 0.00417568
R29425 VDD.n1901 VDD.n635 0.00417568
R29426 VDD.n1513 VDD.n1512 0.00417568
R29427 VDD.n1612 VDD.n1611 0.00417568
R29428 VDD.n1693 VDD.n760 0.00410442
R29429 VDD.n1841 VDD.n1840 0.00410442
R29430 VDD.n443 VDD.n431 0.00408891
R29431 VDD.n453 VDD.n431 0.00408891
R29432 VDD.n454 VDD.n453 0.00408891
R29433 VDD.n455 VDD.n454 0.00408891
R29434 VDD.n465 VDD.n423 0.00408891
R29435 VDD.n466 VDD.n465 0.00408891
R29436 VDD.n467 VDD.n466 0.00408891
R29437 VDD.n467 VDD.n414 0.00408891
R29438 VDD.n478 VDD.n414 0.00408891
R29439 VDD.n479 VDD.n478 0.00408891
R29440 VDD.n480 VDD.n479 0.00408891
R29441 VDD.n480 VDD.n395 0.00408891
R29442 VDD.n550 VDD.n396 0.00408891
R29443 VDD.n546 VDD.n396 0.00408891
R29444 VDD.n546 VDD.n545 0.00408891
R29445 VDD.n545 VDD.n544 0.00408891
R29446 VDD.n544 VDD.n402 0.00408891
R29447 VDD.n510 VDD.n402 0.00408891
R29448 VDD.n511 VDD.n509 0.00408891
R29449 VDD.n515 VDD.n509 0.00408891
R29450 VDD.n516 VDD.n515 0.00408891
R29451 VDD.n517 VDD.n516 0.00408891
R29452 VDD.n517 VDD.n506 0.00408891
R29453 VDD.n521 VDD.n506 0.00408891
R29454 VDD.n1045 VDD.n1037 0.00406757
R29455 VDD.n1254 VDD.n943 0.00406757
R29456 VDD.n1703 VDD.n747 0.00406757
R29457 VDD.n1828 VDD.n1827 0.00406757
R29458 VDD.n831 VDD.n826 0.00402269
R29459 VDD.n1487 VDD.n858 0.00398793
R29460 VDD.n1587 VDD.n802 0.00398793
R29461 VDD.n1317 VDD.n1314 0.00397174
R29462 VDD.n1915 VDD.n1914 0.00397174
R29463 VDD.n1884 VDD.n654 0.00397174
R29464 VDD.n1739 VDD.n1738 0.00394963
R29465 VDD.n1788 VDD.n706 0.00394963
R29466 VDD.n1478 VDD.n871 0.00394626
R29467 VDD.n819 VDD.n814 0.00394626
R29468 VDD.n890 VDD.n872 0.00393696
R29469 VDD.n1560 VDD.n815 0.00393696
R29470 VDD.n862 VDD.n857 0.00390294
R29471 VDD.n1601 VDD.n806 0.00390294
R29472 VDD.n1549 VDD.n827 0.00389381
R29473 VDD.n1507 VDD.n855 0.00385851
R29474 VDD.n1535 VDD.n839 0.00385851
R29475 VDD.n1617 VDD.n1610 0.00385851
R29476 VDD.n789 VDD.n787 0.00385851
R29477 VDD.n1508 VDD.n1507 0.00380768
R29478 VDD.n1617 VDD.n1616 0.00380768
R29479 VDD.n841 VDD.n839 0.00380053
R29480 VDD.n790 VDD.n789 0.00380053
R29481 VDD.n1715 VDD.n742 0.00379484
R29482 VDD.n1816 VDD.n1815 0.00379484
R29483 VDD.n1399 VDD.n953 0.00379484
R29484 VDD.n1675 VDD.n765 0.00377273
R29485 VDD.n1484 VDD.n1483 0.0037725
R29486 VDD.n1549 VDD.n1548 0.0037725
R29487 VDD.n1591 VDD.n1590 0.0037725
R29488 VDD.n1660 VDD.n774 0.00374762
R29489 VDD.n1367 VDD.n1332 0.0037285
R29490 VDD.n1903 VDD.n1902 0.0037285
R29491 VDD.n1362 VDD.n1338 0.00370639
R29492 VDD.n648 VDD.n647 0.00370639
R29493 VDD.n1671 VDD.n1670 0.00369524
R29494 VDD.n1726 VDD.n1725 0.00366216
R29495 VDD.n1807 VDD.n1806 0.00366216
R29496 VDD.n1662 VDD.n777 0.00366216
R29497 VDD.n1657 VDD.n1656 0.00364005
R29498 VDD.n910 VDD.n909 0.00363514
R29499 VDD.n1269 VDD.n945 0.00363514
R29500 VDD.n1697 VDD.n1696 0.00363514
R29501 VDD.n1837 VDD.n1836 0.00363514
R29502 VDD.n1396 VDD.n1395 0.00359048
R29503 VDD.n1544 VDD.n833 0.00358532
R29504 VDD.n1564 VDD.n1561 0.00358218
R29505 VDD.n897 VDD.n896 0.00357902
R29506 VDD.n1292 VDD.n954 0.00357902
R29507 VDD.n1487 VDD.n1486 0.00357098
R29508 VDD.n1588 VDD.n1587 0.00357098
R29509 VDD.n1734 VDD.n1733 0.00348526
R29510 VDD.n1799 VDD.n1798 0.00348526
R29511 VDD.n1511 VDD.n1510 0.003457
R29512 VDD.n1614 VDD.n1613 0.003457
R29513 VDD.n844 VDD.n840 0.00344926
R29514 VDD.n793 VDD.n788 0.00344926
R29515 VDD.n1375 VDD.n1320 0.00344103
R29516 VDD.n1907 VDD.n1906 0.00344103
R29517 VDD.n1889 VDD.n649 0.00344103
R29518 VDD.n1536 VDD.n837 0.00343273
R29519 VDD.n1643 VDD.n1642 0.00343273
R29520 VDD.n1503 VDD.n1502 0.00341839
R29521 VDD.n801 VDD.n800 0.00341839
R29522 VDD.n1608 VDD.n803 0.00341837
R29523 VDD.n1500 VDD.n859 0.00341837
R29524 VDD.n1394 VDD.n1297 0.00335476
R29525 VDD.n1709 VDD.n744 0.00335258
R29526 VDD.n1831 VDD.n1830 0.00335258
R29527 VDD.n1502 VDD.n857 0.0033136
R29528 VDD.n1601 VDD.n801 0.0033136
R29529 VDD.n1005 VDD.n928 0.00331081
R29530 VDD.n1162 VDD.n994 0.00331081
R29531 VDD.n1302 VDD.n1300 0.00331081
R29532 VDD.n1756 VDD.n1755 0.00331081
R29533 VDD.n1776 VDD.n711 0.00331081
R29534 VDD.n1921 VDD.n603 0.00331081
R29535 VDD.n1471 VDD.n870 0.00331081
R29536 VDD.n1579 VDD.n1578 0.00331081
R29537 VDD.n847 VDD.n840 0.00330444
R29538 VDD.n1626 VDD.n788 0.00330444
R29539 VDD.n1539 VDD.n837 0.0032992
R29540 VDD.n1642 VDD.n1641 0.0032992
R29541 VDD.n1510 VDD.n1509 0.00329663
R29542 VDD.n1615 VDD.n1614 0.00329663
R29543 VDD.n1939 VDD.n550 0.00326346
R29544 VDD.n1668 VDD.n775 0.00324201
R29545 VDD.n1753 VDD.n1752 0.00319779
R29546 VDD.n1782 VDD.n708 0.00319779
R29547 VDD.n1866 VDD.n1865 0.00319779
R29548 VDD.n1669 VDD.n773 0.00319779
R29549 VDD.n1391 VDD.n1301 0.00317568
R29550 VDD.n1919 VDD.n1918 0.00317568
R29551 VDD.n1478 VDD.n1477 0.00317568
R29552 VDD.n1585 VDD.n814 0.00317568
R29553 VDD.n1486 VDD.n1485 0.00316007
R29554 VDD.n1589 VDD.n1588 0.00316007
R29555 VDD.n1547 VDD.n833 0.00314581
R29556 VDD.n1296 VDD.n1295 0.00310934
R29557 VDD.n1372 VDD.n1324 0.00309459
R29558 VDD.n633 VDD.n631 0.00309459
R29559 VDD.n1506 VDD.n1505 0.00309459
R29560 VDD.n1619 VDD.n1618 0.00309459
R29561 VDD.n1690 VDD.n1689 0.003043
R29562 VDD.n1855 VDD.n1854 0.003043
R29563 VDD.n1050 VDD.n1048 0.0029881
R29564 VDD.n1085 VDD.n1084 0.0029881
R29565 VDD.n1100 VDD.n1019 0.0029881
R29566 VDD.n1202 VDD.n1201 0.0029881
R29567 VDD.n1485 VDD.n1484 0.00298054
R29568 VDD.n1548 VDD.n1547 0.00298054
R29569 VDD.n1590 VDD.n1589 0.00298054
R29570 VDD.n1217 VDD.n976 0.0029619
R29571 VDD.n1251 VDD.n1250 0.0029619
R29572 VDD.n847 VDD.n841 0.00293083
R29573 VDD.n1626 VDD.n790 0.00293083
R29574 VDD.n1509 VDD.n1508 0.0029237
R29575 VDD.n1616 VDD.n1615 0.0029237
R29576 VDD.n1759 VDD.n719 0.00291032
R29577 VDD.n1763 VDD.n1762 0.00291032
R29578 VDD.n1393 VDD.n1392 0.00291032
R29579 VDD.n606 VDD.n605 0.00291032
R29580 VDD.n1864 VDD.n670 0.00291032
R29581 VDD.n1559 VDD.n826 0.00291032
R29582 VDD.n772 VDD.n771 0.00291032
R29583 VDD.n1503 VDD.n855 0.00289527
R29584 VDD.n1536 VDD.n1535 0.00289527
R29585 VDD.n1610 VDD.n800 0.00289527
R29586 VDD.n1643 VDD.n787 0.00289527
R29587 VDD.n897 VDD.n888 0.00287188
R29588 VDD.n1290 VDD.n954 0.00284569
R29589 VDD.n830 VDD.n827 0.00283826
R29590 VDD.n1859 VDD.n675 0.00283095
R29591 VDD.n875 VDD.n872 0.00279542
R29592 VDD.n818 VDD.n815 0.00279542
R29593 VDD.n861 VDD.n858 0.00276679
R29594 VDD.n805 VDD.n802 0.00276679
R29595 VDD.n755 VDD.n754 0.00275553
R29596 VDD.n1834 VDD.n685 0.00275553
R29597 VDD.n764 VDD.n762 0.00273342
R29598 VDD.n1870 VDD.n671 0.00273342
R29599 VDD.n899 VDD.n888 0.00272619
R29600 VDD.n900 VDD.n899 0.00272619
R29601 VDD.n1459 VDD.n1458 0.00272619
R29602 VDD.n1457 VDD.n906 0.00272619
R29603 VDD.n1448 VDD.n1447 0.00272619
R29604 VDD.n1042 VDD.n1039 0.00272619
R29605 VDD.n1047 VDD.n1039 0.00272619
R29606 VDD.n1049 VDD.n1035 0.00272619
R29607 VDD.n1057 VDD.n1035 0.00272619
R29608 VDD.n1065 VDD.n1032 0.00272619
R29609 VDD.n1066 VDD.n1065 0.00272619
R29610 VDD.n1075 VDD.n1074 0.00272619
R29611 VDD.n1076 VDD.n1075 0.00272619
R29612 VDD.n1086 VDD.n1026 0.00272619
R29613 VDD.n1090 VDD.n1026 0.00272619
R29614 VDD.n1098 VDD.n1022 0.00272619
R29615 VDD.n1099 VDD.n1098 0.00272619
R29616 VDD.n1107 VDD.n1106 0.00272619
R29617 VDD.n1108 VDD.n1016 0.00272619
R29618 VDD.n1120 VDD.n1014 0.00272619
R29619 VDD.n1132 VDD.n1010 0.00272619
R29620 VDD.n1133 VDD.n1132 0.00272619
R29621 VDD.n1139 VDD.n1138 0.00272619
R29622 VDD.n1141 VDD.n1139 0.00272619
R29623 VDD.n1141 VDD.n1140 0.00272619
R29624 VDD.n1150 VDD.n1149 0.00272619
R29625 VDD.n1159 VDD.n1158 0.00272619
R29626 VDD.n1158 VDD.n996 0.00272619
R29627 VDD.n1168 VDD.n1167 0.00272619
R29628 VDD.n1167 VDD.n992 0.00272619
R29629 VDD.n1174 VDD.n992 0.00272619
R29630 VDD.n1182 VDD.n989 0.00272619
R29631 VDD.n1183 VDD.n1182 0.00272619
R29632 VDD.n1192 VDD.n1191 0.00272619
R29633 VDD.n1193 VDD.n1192 0.00272619
R29634 VDD.n1207 VDD.n983 0.00272619
R29635 VDD.n1216 VDD.n1215 0.00272619
R29636 VDD.n1224 VDD.n1223 0.00272619
R29637 VDD.n1225 VDD.n973 0.00272619
R29638 VDD.n1237 VDD.n971 0.00272619
R29639 VDD.n1249 VDD.n967 0.00272619
R29640 VDD.n1250 VDD.n1249 0.00272619
R29641 VDD.n1257 VDD.n965 0.00272619
R29642 VDD.n1258 VDD.n1257 0.00272619
R29643 VDD.n1259 VDD.n1258 0.00272619
R29644 VDD.n1266 VDD.n1265 0.00272619
R29645 VDD.n1266 VDD.n959 0.00272619
R29646 VDD.n1274 VDD.n957 0.00272619
R29647 VDD.n1281 VDD.n957 0.00272619
R29648 VDD.n1288 VDD.n1287 0.00272619
R29649 VDD.n1290 VDD.n1289 0.00272619
R29650 VDD.n900 VDD.n885 0.0027
R29651 VDD.n1458 VDD.n1457 0.0027
R29652 VDD.n1448 VDD.n908 0.0027
R29653 VDD.n1042 VDD.n1041 0.0027
R29654 VDD.n1050 VDD.n1049 0.0027
R29655 VDD.n1076 VDD.n1028 0.0027
R29656 VDD.n1108 VDD.n1107 0.0027
R29657 VDD.n1116 VDD.n1014 0.0027
R29658 VDD.n1122 VDD.n1010 0.0027
R29659 VDD.n1150 VDD.n1148 0.0027
R29660 VDD.n1159 VDD.n1157 0.0027
R29661 VDD.n1193 VDD.n985 0.0027
R29662 VDD.n1203 VDD.n983 0.0027
R29663 VDD.n1215 VDD.n979 0.0027
R29664 VDD.n1225 VDD.n1224 0.0027
R29665 VDD.n1233 VDD.n971 0.0027
R29666 VDD.n1239 VDD.n967 0.0027
R29667 VDD.n1282 VDD.n1281 0.0027
R29668 VDD.n1289 VDD.n1288 0.0027
R29669 VDD.n1084 VDD.n1028 0.00264762
R29670 VDD.n1223 VDD.n976 0.00264762
R29671 VDD.n1378 VDD.n1315 0.00264496
R29672 VDD.n626 VDD.n625 0.00264496
R29673 VDD.n1888 VDD.n652 0.00262285
R29674 VDD.n1540 VDD.n835 0.00262285
R29675 VDD.n1640 VDD.n1637 0.00262285
R29676 VDD.n1100 VDD.n1099 0.00262143
R29677 VDD.n1203 VDD.n1202 0.00262143
R29678 VDD.n732 VDD.n729 0.00260074
R29679 VDD.n1786 VDD.n698 0.00260074
R29680 VDD.n1052 VDD.n1038 0.00257862
R29681 VDD.n1252 VDD.n966 0.00257862
R29682 VDD.n1201 VDD.n985 0.00256905
R29683 VDD.n1096 VDD.n923 0.00255405
R29684 VDD.n1197 VDD.n981 0.00255405
R29685 VDD.n1731 VDD.n1730 0.00255405
R29686 VDD.n1796 VDD.n697 0.00255405
R29687 VDD.n1106 VDD.n1019 0.00254286
R29688 VDD.n1217 VDD.n1216 0.00254286
R29689 VDD.n1102 VDD.n1020 0.0025344
R29690 VDD.n1086 VDD.n1085 0.00251667
R29691 VDD.n1200 VDD.n1199 0.00251228
R29692 VDD.n1565 VDD.n1564 0.00249519
R29693 VDD.n894 VDD.n893 0.0024936
R29694 VDD.n1048 VDD.n1047 0.00246429
R29695 VDD.n1251 VDD.n965 0.00246429
R29696 VDD.n1713 VDD.n734 0.00244595
R29697 VDD.n1810 VDD.n694 0.00244595
R29698 VDD.n1067 VDD.n1066 0.0024381
R29699 VDD.n1233 VDD.n1232 0.0024381
R29700 VDD.n1083 VDD.n1082 0.00242383
R29701 VDD.n1219 VDD.n977 0.00242383
R29702 VDD.n1661 VDD.n1660 0.00238571
R29703 VDD.n1397 VDD.n1396 0.00238571
R29704 VDD.n1453 VDD.n1452 0.00238571
R29705 VDD.n1446 VDD.n913 0.00238571
R29706 VDD.n1059 VDD.n1058 0.00238571
R29707 VDD.n1067 VDD.n1030 0.00238571
R29708 VDD.n1092 VDD.n1091 0.00238571
R29709 VDD.n1115 VDD.n1114 0.00238571
R29710 VDD.n1123 VDD.n1121 0.00238571
R29711 VDD.n1147 VDD.n1003 0.00238571
R29712 VDD.n1156 VDD.n999 0.00238571
R29713 VDD.n1165 VDD.n996 0.00238571
R29714 VDD.n1176 VDD.n1175 0.00238571
R29715 VDD.n1184 VDD.n987 0.00238571
R29716 VDD.n1209 VDD.n1208 0.00238571
R29717 VDD.n1232 VDD.n1231 0.00238571
R29718 VDD.n1240 VDD.n1238 0.00238571
R29719 VDD.n1264 VDD.n963 0.00238571
R29720 VDD.n1273 VDD.n1272 0.00238571
R29721 VDD.n1460 VDD.n884 0.00237961
R29722 VDD.n1456 VDD.n1455 0.00237961
R29723 VDD.n1449 VDD.n912 0.00237961
R29724 VDD.n1044 VDD.n1043 0.00237961
R29725 VDD.n1046 VDD.n1044 0.00237961
R29726 VDD.n1055 VDD.n1036 0.00237961
R29727 VDD.n1056 VDD.n1055 0.00237961
R29728 VDD.n1064 VDD.n1033 0.00237961
R29729 VDD.n1064 VDD.n1031 0.00237961
R29730 VDD.n1073 VDD.n1029 0.00237961
R29731 VDD.n1077 VDD.n1029 0.00237961
R29732 VDD.n1088 VDD.n1087 0.00237961
R29733 VDD.n1089 VDD.n1088 0.00237961
R29734 VDD.n1097 VDD.n1023 0.00237961
R29735 VDD.n1097 VDD.n1021 0.00237961
R29736 VDD.n1105 VDD.n1018 0.00237961
R29737 VDD.n1109 VDD.n1017 0.00237961
R29738 VDD.n1119 VDD.n1118 0.00237961
R29739 VDD.n1131 VDD.n1130 0.00237961
R29740 VDD.n1131 VDD.n1009 0.00237961
R29741 VDD.n1137 VDD.n1006 0.00237961
R29742 VDD.n1142 VDD.n1006 0.00237961
R29743 VDD.n1142 VDD.n1007 0.00237961
R29744 VDD.n1151 VDD.n1002 0.00237961
R29745 VDD.n1160 VDD.n997 0.00237961
R29746 VDD.n1163 VDD.n997 0.00237961
R29747 VDD.n1169 VDD.n993 0.00237961
R29748 VDD.n1172 VDD.n993 0.00237961
R29749 VDD.n1173 VDD.n1172 0.00237961
R29750 VDD.n1181 VDD.n990 0.00237961
R29751 VDD.n1181 VDD.n988 0.00237961
R29752 VDD.n1190 VDD.n986 0.00237961
R29753 VDD.n1194 VDD.n986 0.00237961
R29754 VDD.n1206 VDD.n1205 0.00237961
R29755 VDD.n1214 VDD.n978 0.00237961
R29756 VDD.n1222 VDD.n975 0.00237961
R29757 VDD.n1226 VDD.n974 0.00237961
R29758 VDD.n1236 VDD.n1235 0.00237961
R29759 VDD.n1248 VDD.n1247 0.00237961
R29760 VDD.n1248 VDD.n966 0.00237961
R29761 VDD.n1256 VDD.n1255 0.00237961
R29762 VDD.n1256 VDD.n964 0.00237961
R29763 VDD.n1260 VDD.n964 0.00237961
R29764 VDD.n1267 VDD.n962 0.00237961
R29765 VDD.n1267 VDD.n960 0.00237961
R29766 VDD.n1279 VDD.n1275 0.00237961
R29767 VDD.n1280 VDD.n1279 0.00237961
R29768 VDD.n1286 VDD.n951 0.00237961
R29769 VDD.n1366 VDD.n1365 0.00237961
R29770 VDD.n1365 VDD.n1333 0.00237961
R29771 VDD.n645 VDD.n630 0.00237961
R29772 VDD.n646 VDD.n645 0.00237961
R29773 VDD.n892 VDD.n887 0.00237961
R29774 VDD.n1473 VDD.n1472 0.00237961
R29775 VDD.n1530 VDD.n843 0.00237961
R29776 VDD.n1530 VDD.n1529 0.00237961
R29777 VDD.n1555 VDD.n1554 0.00237961
R29778 VDD.n1581 VDD.n1580 0.00237961
R29779 VDD.n1632 VDD.n792 0.00237961
R29780 VDD.n1632 VDD.n1631 0.00237961
R29781 VDD.n1116 VDD.n1115 0.00235952
R29782 VDD.n1138 VDD.n1008 0.00235952
R29783 VDD.n902 VDD.n901 0.00235749
R29784 VDD.n1456 VDD.n884 0.00235749
R29785 VDD.n1450 VDD.n1449 0.00235749
R29786 VDD.n1043 VDD.n1040 0.00235749
R29787 VDD.n1051 VDD.n1036 0.00235749
R29788 VDD.n1078 VDD.n1077 0.00235749
R29789 VDD.n1109 VDD.n1018 0.00235749
R29790 VDD.n1118 VDD.n1117 0.00235749
R29791 VDD.n1130 VDD.n1011 0.00235749
R29792 VDD.n1151 VDD.n1001 0.00235749
R29793 VDD.n1160 VDD.n998 0.00235749
R29794 VDD.n1195 VDD.n1194 0.00235749
R29795 VDD.n1205 VDD.n1204 0.00235749
R29796 VDD.n1214 VDD.n980 0.00235749
R29797 VDD.n1226 VDD.n975 0.00235749
R29798 VDD.n1235 VDD.n1234 0.00235749
R29799 VDD.n1247 VDD.n968 0.00235749
R29800 VDD.n1280 VDD.n956 0.00235749
R29801 VDD.n1498 VDD.n1497 0.00235749
R29802 VDD.n1606 VDD.n1605 0.00235749
R29803 VDD.n1184 VDD.n1183 0.00233333
R29804 VDD.n1083 VDD.n1078 0.00231327
R29805 VDD.n1222 VDD.n977 0.00231327
R29806 VDD.n904 VDD.n885 0.00230714
R29807 VDD.n1283 VDD.n1282 0.00230714
R29808 VDD.n1287 VDD.n955 0.00230714
R29809 VDD.n1101 VDD.n1021 0.00229115
R29810 VDD.n1204 VDD.n984 0.00229115
R29811 VDD.n1714 VDD.n1713 0.00229115
R29812 VDD.n1817 VDD.n1810 0.00229115
R29813 VDD.n1459 VDD.n905 0.00228095
R29814 VDD.n1447 VDD.n1446 0.00228095
R29815 VDD.n1265 VDD.n1264 0.00225476
R29816 VDD.n1200 VDD.n1195 0.00224693
R29817 VDD.n1389 VDD.n1303 0.00222973
R29818 VDD.n611 VDD.n604 0.00222973
R29819 VDD.n1481 VDD.n1480 0.00222973
R29820 VDD.n1593 VDD.n811 0.00222973
R29821 VDD.n1105 VDD.n1020 0.00222482
R29822 VDD.n1218 VDD.n978 0.00222482
R29823 VDD.n1087 VDD.n1027 0.0022027
R29824 VDD.n1134 VDD.n1133 0.00220238
R29825 VDD.n1168 VDD.n1166 0.00220238
R29826 VDD.n1148 VDD.n1147 0.00217619
R29827 VDD.n1149 VDD.n999 0.00217619
R29828 VDD.n1561 VDD.n1560 0.00217613
R29829 VDD.n1046 VDD.n1038 0.00215848
R29830 VDD.n1255 VDD.n1252 0.00215848
R29831 VDD.n1068 VDD.n1031 0.00213636
R29832 VDD.n1234 VDD.n972 0.00213636
R29833 VDD.n1740 VDD.n729 0.00213636
R29834 VDD.n1787 VDD.n1786 0.00213636
R29835 VDD.n1885 VDD.n652 0.00211425
R29836 VDD.n1543 VDD.n835 0.00211425
R29837 VDD.n1637 VDD.n779 0.00211425
R29838 VDD.n1395 VDD.n1394 0.00209762
R29839 VDD.n1452 VDD.n908 0.00209762
R29840 VDD.n1164 VDD.n1163 0.00209214
R29841 VDD.n1379 VDD.n1378 0.00209214
R29842 VDD.n625 VDD.n610 0.00209214
R29843 VDD.n1499 VDD.n861 0.00209214
R29844 VDD.n1607 VDD.n805 0.00209214
R29845 VDD.n1272 VDD.n959 0.00207143
R29846 VDD.n1117 VDD.n1015 0.00207002
R29847 VDD.n1137 VDD.n1136 0.00207002
R29848 VDD.n1185 VDD.n988 0.00204791
R29849 VDD.n903 VDD.n902 0.0020258
R29850 VDD.n1284 VDD.n956 0.0020258
R29851 VDD.n1286 VDD.n1285 0.0020258
R29852 VDD.n1121 VDD.n1120 0.00201905
R29853 VDD.n1323 VDD.n1322 0.00201351
R29854 VDD.n1909 VDD.n1908 0.00201351
R29855 VDD.n1495 VDD.n856 0.00201351
R29856 VDD.n1603 VDD.n1602 0.00201351
R29857 VDD.n1460 VDD.n883 0.00200369
R29858 VDD.n1445 VDD.n912 0.00200369
R29859 VDD.n756 VDD.n755 0.00200369
R29860 VDD.n1835 VDD.n1834 0.00200369
R29861 VDD.n1398 VDD.n1293 0.00200107
R29862 VDD.n895 VDD.n894 0.00200107
R29863 VDD.n893 VDD.n874 0.00200107
R29864 VDD.n1176 VDD.n989 0.00199286
R29865 VDD.n1263 VDD.n962 0.00198157
R29866 VDD.n1135 VDD.n1009 0.00193735
R29867 VDD.n1169 VDD.n995 0.00193735
R29868 VDD.n1146 VDD.n1001 0.00191523
R29869 VDD.n1002 VDD.n1000 0.00191523
R29870 VDD.n1399 VDD.n952 0.00191523
R29871 VDD.n1870 VDD.n674 0.00191523
R29872 VDD.n898 VDD.n887 0.00191523
R29873 VDD.n892 VDD.n891 0.00191523
R29874 VDD.n1059 VDD.n1032 0.00191429
R29875 VDD.n1238 VDD.n1237 0.00191429
R29876 VDD.n1072 VDD.n1071 0.00187101
R29877 VDD.n1497 VDD.n862 0.00185493
R29878 VDD.n1605 VDD.n806 0.00185493
R29879 VDD.n1451 VDD.n1450 0.00184889
R29880 VDD.n1230 VDD.n1229 0.00184889
R29881 VDD.n1759 VDD.n1758 0.00184889
R29882 VDD.n1766 VDD.n1763 0.00184889
R29883 VDD.n1393 VDD.n1296 0.00184889
R29884 VDD.n605 VDD.n597 0.00184889
R29885 VDD.n1872 VDD.n670 0.00184889
R29886 VDD.n1474 VDD.n875 0.00184889
R29887 VDD.n1567 VDD.n1559 0.00184889
R29888 VDD.n1582 VDD.n818 0.00184889
R29889 VDD.n1677 VDD.n771 0.00184889
R29890 VDD.n1209 VDD.n979 0.00183571
R29891 VDD.n1271 VDD.n960 0.00182678
R29892 VDD.n1091 VDD.n1090 0.00180952
R29893 VDD.n1080 VDD.n1024 0.0017973
R29894 VDD.n1213 VDD.n938 0.0017973
R29895 VDD.n1723 VDD.n733 0.0017973
R29896 VDD.n1804 VDD.n1803 0.0017973
R29897 VDD.n1472 VDD.n871 0.0017897
R29898 VDD.n1580 VDD.n819 0.0017897
R29899 VDD.n1113 VDD.n1112 0.00178256
R29900 VDD.n1119 VDD.n1013 0.00178256
R29901 VDD.n1189 VDD.n1188 0.00178256
R29902 VDD.n1177 VDD.n990 0.00176044
R29903 VDD.n1670 VDD.n774 0.00175714
R29904 VDD.n1092 VDD.n1022 0.00173095
R29905 VDD.n1208 VDD.n1207 0.00173095
R29906 VDD.n1444 VDD.n914 0.00171622
R29907 VDD.n1554 VDD.n831 0.00171347
R29908 VDD.n1060 VDD.n1033 0.0016941
R29909 VDD.n1236 VDD.n970 0.0016941
R29910 VDD.n1262 VDD.n1261 0.0016941
R29911 VDD.n1690 VDD.n753 0.0016941
R29912 VDD.n1855 VDD.n677 0.0016941
R29913 VDD.n1240 VDD.n1239 0.00165238
R29914 VDD.n1145 VDD.n1004 0.00162776
R29915 VDD.n1155 VDD.n1154 0.00162776
R29916 VDD.n1210 VDD.n980 0.00162776
R29917 VDD.n1295 VDD.n1294 0.00162776
R29918 VDD.n1058 VDD.n1057 0.00162619
R29919 VDD.n1089 VDD.n1025 0.00160565
R29920 VDD.n1388 VDD.n1301 0.00158354
R29921 VDD.n1918 VDD.n607 0.00158354
R29922 VDD.n1477 VDD.n869 0.00158354
R29923 VDD.n1586 VDD.n1585 0.00158354
R29924 VDD.n1454 VDD.n907 0.00156143
R29925 VDD.n1270 VDD.n958 0.00156143
R29926 VDD.n1752 VDD.n1751 0.00156143
R29927 VDD.n1782 VDD.n1781 0.00156143
R29928 VDD.n1866 VDD.n656 0.00156143
R29929 VDD.n1556 VDD.n830 0.00156143
R29930 VDD.n1669 VDD.n1668 0.00156143
R29931 VDD.n1123 VDD.n1122 0.00154762
R29932 VDD.n1175 VDD.n1174 0.00154762
R29933 VDD.n1093 VDD.n1023 0.00153931
R29934 VDD.n1206 VDD.n982 0.00153931
R29935 VDD.n1125 VDD.n1124 0.00149509
R29936 VDD.n1663 VDD.n775 0.00149509
R29937 VDD.n1178 VDD.n991 0.00147297
R29938 VDD.n1241 VDD.n968 0.00147297
R29939 VDD.n1453 VDD.n906 0.00146905
R29940 VDD.n1274 VDD.n1273 0.00146905
R29941 VDD.n1056 VDD.n1034 0.00145086
R29942 VDD.n1061 VDD.n1034 0.00140663
R29943 VDD.n1242 VDD.n1241 0.00140663
R29944 VDD.n1709 VDD.n1708 0.00140663
R29945 VDD.n1831 VDD.n687 0.00140663
R29946 VDD.n1157 VDD.n1156 0.00139048
R29947 VDD.n1124 VDD.n1011 0.00138452
R29948 VDD.n1173 VDD.n991 0.00138452
R29949 VDD.n905 VDD.n904 0.00136429
R29950 VDD.n1134 VDD.n1008 0.00136429
R29951 VDD.n1140 VDD.n1003 0.00136429
R29952 VDD.n1094 VDD.n1093 0.00134029
R29953 VDD.n1211 VDD.n982 0.00134029
R29954 VDD.n1166 VDD.n1165 0.00133809
R29955 VDD.n1283 VDD.n955 0.00133809
R29956 VDD.n1939 VDD.n395 0.00132545
R29957 VDD.n1455 VDD.n1454 0.00131818
R29958 VDD.n1275 VDD.n958 0.00131818
R29959 VDD.n1556 VDD.n1555 0.00131818
R29960 VDD.n1375 VDD.n1374 0.00129607
R29961 VDD.n1336 VDD.n587 0.00129607
R29962 VDD.n1906 VDD.n627 0.00129607
R29963 VDD.n1892 VDD.n649 0.00129607
R29964 VDD.n1041 VDD.n913 0.00128571
R29965 VDD.n1259 VDD.n963 0.00128571
R29966 VDD.n1094 VDD.n1025 0.00125184
R29967 VDD.n1155 VDD.n998 0.00125184
R29968 VDD.n1211 VDD.n1210 0.00125184
R29969 VDD.n1734 VDD.n731 0.00125184
R29970 VDD.n1800 VDD.n1799 0.00125184
R29971 VDD.n903 VDD.n883 0.00122973
R29972 VDD.n1136 VDD.n1135 0.00122973
R29973 VDD.n1007 VDD.n1004 0.00122973
R29974 VDD.n1164 VDD.n995 0.00120762
R29975 VDD.n1285 VDD.n1284 0.00120762
R29976 VDD.n1114 VDD.n1016 0.00120714
R29977 VDD.n1191 VDD.n987 0.00120714
R29978 VDD.n1061 VDD.n1060 0.0011855
R29979 VDD.n1242 VDD.n970 0.0011855
R29980 VDD.n1040 VDD.n914 0.00116339
R29981 VDD.n1261 VDD.n1260 0.00116339
R29982 VDD.n1385 VDD.n1384 0.00114865
R29983 VDD.n615 VDD.n614 0.00114865
R29984 VDD.n1489 VDD.n867 0.00114865
R29985 VDD.n813 VDD.n812 0.00114865
R29986 VDD.n1231 VDD.n973 0.00112857
R29987 VDD.n1178 VDD.n1177 0.00111916
R29988 VDD.n1074 VDD.n1030 0.00110238
R29989 VDD.n1113 VDD.n1017 0.00109705
R29990 VDD.n1125 VDD.n1013 0.00109705
R29991 VDD.n1190 VDD.n1189 0.00109705
R29992 VDD.n1727 VDD.n1726 0.00109705
R29993 VDD.n1807 VDD.n696 0.00109705
R29994 VDD.n1663 VDD.n1662 0.00109705
R29995 VDD.n1362 VDD.n1361 0.00105283
R29996 VDD.n1894 VDD.n648 0.00105283
R29997 VDD.n1858 VDD.n674 0.00105283
R29998 VDD.n1144 VDD.n929 0.00104054
R29999 VDD.n1770 VDD.n715 0.00104054
R30000 VDD.n1451 VDD.n907 0.00103071
R30001 VDD.n1230 VDD.n974 0.00103071
R30002 VDD.n1271 VDD.n1270 0.00103071
R30003 VDD.n1291 VDD.n952 0.00103071
R30004 VDD.n1332 VDD.n1331 0.00103071
R30005 VDD.n1903 VDD.n629 0.00103071
R30006 VDD.n898 VDD.n889 0.00103071
R30007 VDD.n1474 VDD.n1473 0.00103071
R30008 VDD.n1582 VDD.n1581 0.00103071
R30009 VDD.n581 VDD.n578 0.00102022
R30010 VDD.n1073 VDD.n1072 0.0010086
R30011 VDD.n1146 VDD.n1145 0.000964373
R30012 VDD.n1154 VDD.n1000 0.000964373
R30013 VDD.n1294 VDD.n953 0.000964373
R30014 VDD.n891 VDD.n890 0.000964373
R30015 VDD.n1676 VDD.n1675 0.000964373
R30016 VDD.n745 VDD.n742 0.00094226
R30017 VDD.n1815 VDD.n1814 0.00094226
R30018 VDD.n1381 VDD.n1380 0.000932432
R30019 VDD.n1912 VDD.n616 0.000932432
R30020 VDD.n868 VDD.n863 0.000932432
R30021 VDD.n1600 VDD.n1599 0.000932432
R30022 VDD.n901 VDD.n887 0.000898034
R30023 VDD.n1263 VDD.n1262 0.000898034
R30024 VDD.n1445 VDD.n1444 0.000875921
R30025 VDD.n1399 VDD.n951 0.000853808
R30026 VDD.n1656 VDD.n1655 0.000831695
R30027 VDD.n1659 VDD.n1658 0.000814286
R30028 VDD.n1112 VDD.n1015 0.000809582
R30029 VDD.n1188 VDD.n1185 0.000809582
R30030 VDD.n1738 VDD.n721 0.000787469
R30031 VDD.n709 VDD.n706 0.000787469
R30032 VDD.n1499 VDD.n1498 0.000787469
R30033 VDD.n1607 VDD.n1606 0.000787469
R30034 VDD.n1317 VDD.n1304 0.000765356
R30035 VDD.n1915 VDD.n609 0.000765356
R30036 VDD.n1881 VDD.n654 0.000765356
R30037 VDD.n1657 VDD.n777 0.000765356
R30038 VDD.n1229 VDD.n972 0.000743243
R30039 VDD.n1071 VDD.n1068 0.00072113
R30040 VDD.n1443 VDD.n1442 0.000716216
R30041 VDD.n961 VDD.n944 0.000716216
R30042 VDD.n759 VDD.n758 0.000716216
R30043 VDD.n1843 VDD.n1842 0.000716216
R30044 VDD.n1082 VDD.n1027 0.000676904
R30045 VDD.n1219 VDD.n1218 0.000654791
R30046 VDD.n1694 VDD.n1693 0.000654791
R30047 VDD.n1840 VDD.n1839 0.000654791
R30048 VDD.n1199 VDD.n984 0.000588452
R30049 VDD.n1102 VDD.n1101 0.000566339
R30050 VDD.n1052 VDD.n1051 0.000522113
R30051 VDD.n765 VDD.n764 0.000522113
C1083 Y2 VSS 0.12039p
C1084 X2 VSS 91.68561f
C1085 Y1 VSS 0.10102p
C1086 X1 VSS 94.7177f
C1087 CLK_OUT VSS 92.2343f
C1088 Y0 VSS 92.142f
C1089 X0 VSS 90.2415f
C1090 CLK_IN VSS 93.6639f
C1091 nEN VSS 0.10244p
C1092 VDD VSS 0.19687p
C1093 m7_16847_2260# VSS 93.0612f
C1094 m6_60810_42209# VSS 1.80367f
C1095 m6_17427_2840# VSS 0.10708p
C1096 m6_16847_2260# VSS 0.11472p
C1097 m5_17331_2744# VSS 79.2024f
C1098 m5_16847_2260# VSS 84.4749f
C1099 m4_17285_2698# VSS 84.41901f
C1100 m4_16847_2260# VSS 89.24989f
C1101 m3_17285_2698# VSS 91.8291f
C1102 m3_16847_2260# VSS 96.21301f
C1103 m2_17285_2698# VSS 0.10557p
C1104 m2_16847_2260# VSS 0.10679p
C1105 m1_17285_2698# VSS 0.22685p
C1106 m1_16847_2260# VSS 0.22893p
C1107 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.nQ VSS 0.08893f $ **FLOATING
C1108 a_62900_20179# VSS 0.34783f $ **FLOATING
C1109 a_63463_20216# VSS 0.43565f $ **FLOATING
C1110 a_62654_20215# VSS 0.80634f $ **FLOATING
C1111 a_62119_20605# VSS 0.26895f $ **FLOATING
C1112 a_62270_20543# VSS 0.16883f $ **FLOATING
C1113 a_61887_20534# VSS 1.05953f $ **FLOATING
C1114 a_61394_20220# VSS 0.13262f $ **FLOATING
C1115 a_61691_20534# VSS 0.79964f $ **FLOATING
C1116 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.sg13g2_dfrbp_1_0.CLK VSS 0.51487f $ **FLOATING
C1117 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.sg13g2_dfrbp_1_0.CLK VSS 0.51489f $ **FLOATING
C1118 a_54504_20259# VSS 0.13262f $ **FLOATING
C1119 a_53899_20488# VSS 0.16883f $ **FLOATING
C1120 a_53968_20434# VSS 0.26896f $ **FLOATING
C1121 a_53738_20514# VSS 1.05953f $ **FLOATING
C1122 a_53445_20214# VSS 0.34783f $ **FLOATING
C1123 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.nQ VSS 0.08893f $ **FLOATING
C1124 a_53774_20178# VSS 0.80054f $ **FLOATING
C1125 a_53065_20179# VSS 0.80634f $ **FLOATING
C1126 a_52950_20401# VSS 0.43566f $ **FLOATING
C1127 a_64384_21091# VSS 0.59054f $ **FLOATING
C1128 3bit_freq_divider_1.sg13g2_or3_1_0.A VSS 0.77543f $ **FLOATING
C1129 a_63255_21488# VSS 0.38381f $ **FLOATING
C1130 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.D VSS 0.49782f $ **FLOATING
C1131 a_61707_21488# VSS 0.36496f $ **FLOATING
C1132 3bit_freq_divider_1.freq_div_cell_1.Cout VSS 0.14556f $ **FLOATING
C1133 a_60967_21478# VSS 0.27989f $ **FLOATING
C1134 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.Q VSS 2.25165f $ **FLOATING
C1135 3bit_freq_divider_0.freq_div_cell_1.Cout VSS 0.14556f $ **FLOATING
C1136 a_55345_21385# VSS 0.27989f $ **FLOATING
C1137 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.D VSS 0.49784f $ **FLOATING
C1138 a_54434_21392# VSS 0.36496f $ **FLOATING
C1139 3bit_freq_divider_0.sg13g2_or3_1_0.A VSS 0.77447f $ **FLOATING
C1140 a_51648_21103# VSS 0.59026f $ **FLOATING
C1141 a_52886_21392# VSS 0.3838f $ **FLOATING
C1142 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.Q VSS 2.25169f $ **FLOATING
C1143 a_60922_21796# VSS 0.03012f $ **FLOATING
C1144 a_60922_21818# VSS 0.02768f $ **FLOATING
C1145 a_52808_21795# VSS 0.03012f $ **FLOATING
C1146 a_52808_21817# VSS 0.02768f $ **FLOATING
C1147 3bit_freq_divider_1.dff_nclk_0.sg13g2_dfrbp_1_0.CLK VSS 0.50854f $ **FLOATING
C1148 a_64424_22200# VSS 0.12168f $ **FLOATING
C1149 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.nQ VSS 0.07921f $ **FLOATING
C1150 a_62900_21935# VSS 0.33549f $ **FLOATING
C1151 a_63463_21972# VSS 0.42316f $ **FLOATING
C1152 a_62654_21971# VSS 0.7639f $ **FLOATING
C1153 a_62119_22361# VSS 0.25006f $ **FLOATING
C1154 a_62270_22299# VSS 0.1501f $ **FLOATING
C1155 a_61887_22290# VSS 1.02135f $ **FLOATING
C1156 a_61394_21976# VSS 0.12168f $ **FLOATING
C1157 a_61691_22290# VSS 0.77938f $ **FLOATING
C1158 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK VSS 0.47143f $ **FLOATING
C1159 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK VSS 0.47143f $ **FLOATING
C1160 a_54504_22015# VSS 0.12168f $ **FLOATING
C1161 a_53899_22244# VSS 0.1501f $ **FLOATING
C1162 a_53968_22190# VSS 0.25006f $ **FLOATING
C1163 a_53738_22270# VSS 1.02135f $ **FLOATING
C1164 a_53445_21970# VSS 0.33549f $ **FLOATING
C1165 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.nQ VSS 0.07921f $ **FLOATING
C1166 a_53774_21934# VSS 0.78026f $ **FLOATING
C1167 a_53065_21935# VSS 0.7639f $ **FLOATING
C1168 a_52950_22157# VSS 0.4233f $ **FLOATING
C1169 3bit_freq_divider_1.sg13g2_or3_1_0.B VSS 1.39257f $ **FLOATING
C1170 a_64383_23300# VSS 0.25093f $ **FLOATING
C1171 a_63255_23244# VSS 0.37914f $ **FLOATING
C1172 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.D VSS 0.45601f $ **FLOATING
C1173 a_61707_23244# VSS 0.36159f $ **FLOATING
C1174 3bit_freq_divider_1.freq_div_cell_0.Cout VSS 1.80113f $ **FLOATING
C1175 a_60967_23234# VSS 0.27786f $ **FLOATING
C1176 a_64419_23326# VSS 0.1501f $ **FLOATING
C1177 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.Q VSS 2.24178f $ **FLOATING
C1178 3bit_freq_divider_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK VSS 0.50854f $ **FLOATING
C1179 a_51684_22284# VSS 0.12168f $ **FLOATING
C1180 3bit_freq_divider_0.freq_div_cell_0.Cout VSS 1.80115f $ **FLOATING
C1181 a_55345_23141# VSS 0.27786f $ **FLOATING
C1182 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.D VSS 0.45601f $ **FLOATING
C1183 a_54434_23148# VSS 0.36159f $ **FLOATING
C1184 3bit_freq_divider_0.sg13g2_or3_1_0.B VSS 1.39146f $ **FLOATING
C1185 a_52886_23148# VSS 0.37912f $ **FLOATING
C1186 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.Q VSS 2.2418f $ **FLOATING
C1187 a_64383_23628# VSS 0.82074f $ **FLOATING
C1188 a_64383_23434# VSS 1.02665f $ **FLOATING
C1189 a_60922_23552# VSS 0.03012f $ **FLOATING
C1190 a_60922_23574# VSS 0.02768f $ **FLOATING
C1191 a_52808_23551# VSS 0.03012f $ **FLOATING
C1192 a_52808_23573# VSS 0.02768f $ **FLOATING
C1193 a_51693_23426# VSS 0.25093f $ **FLOATING
C1194 a_51693_23075# VSS 0.1501f $ **FLOATING
C1195 a_64383_23706# VSS 0.33666f $ **FLOATING
C1196 3bit_freq_divider_1.dff_nclk_0.D VSS 0.57206f $ **FLOATING
C1197 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.nQ VSS 0.08281f $ **FLOATING
C1198 a_62900_23691# VSS 0.33612f $ **FLOATING
C1199 a_63463_23728# VSS 0.42235f $ **FLOATING
C1200 a_62654_23727# VSS 0.76426f $ **FLOATING
C1201 a_62119_24117# VSS 0.25006f $ **FLOATING
C1202 a_62270_24055# VSS 0.1501f $ **FLOATING
C1203 a_61887_24046# VSS 1.02191f $ **FLOATING
C1204 a_61394_23732# VSS 0.12168f $ **FLOATING
C1205 a_61691_24046# VSS 0.78738f $ **FLOATING
C1206 3bit_freq_divider_1.dff_nclk_0.nCLK VSS 7.48134f $ **FLOATING
C1207 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.sg13g2_dfrbp_1_0.CLK VSS 0.47246f $ **FLOATING
C1208 a_51631_22774# VSS 0.82147f $ **FLOATING
C1209 a_51684_22692# VSS 1.02713f $ **FLOATING
C1210 3bit_freq_divider_1.sg13g2_nand2_1_0.Y VSS 2.56526f $ **FLOATING
C1211 3bit_freq_divider_0.sg13g2_nand2_1_0.Y VSS 2.56527f $ **FLOATING
C1212 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.sg13g2_dfrbp_1_0.CLK VSS 0.47246f $ **FLOATING
C1213 a_54504_23771# VSS 0.12168f $ **FLOATING
C1214 a_53899_24000# VSS 0.1501f $ **FLOATING
C1215 a_53968_23946# VSS 0.25006f $ **FLOATING
C1216 a_53738_24026# VSS 1.02191f $ **FLOATING
C1217 a_53445_23726# VSS 0.33612f $ **FLOATING
C1218 3bit_freq_divider_0.dff_nclk_0.nCLK VSS 7.50548f $ **FLOATING
C1219 a_51685_23725# VSS 0.33666f $ **FLOATING
C1220 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.nQ VSS 0.08281f $ **FLOATING
C1221 a_53774_23690# VSS 0.78853f $ **FLOATING
C1222 a_53065_23691# VSS 0.76426f $ **FLOATING
C1223 a_52950_23913# VSS 0.42231f $ **FLOATING
C1224 a_64383_23889# VSS 0.79267f $ **FLOATING
C1225 a_64384_24445# VSS 0.41218f $ **FLOATING
C1226 3bit_freq_divider_0.dff_nclk_0.D VSS 0.57206f $ **FLOATING
C1227 a_51648_24041# VSS 0.7928f $ **FLOATING
C1228 3bit_freq_divider_1.dff_nclk_0.nRST VSS 1.21235f $ **FLOATING
C1229 a_64398_24796# VSS 0.17085f $ **FLOATING
C1230 a_64338_24910# VSS 0.01158f $ **FLOATING
C1231 a_64362_24865# VSS 0.18902f $ **FLOATING
C1232 a_64459_24995# VSS 0.21807f $ **FLOATING
C1233 a_51648_24438# VSS 0.41218f $ **FLOATING
C1234 3bit_freq_divider_1.sg13g2_or3_1_0.C VSS 2.00849f $ **FLOATING
C1235 a_63255_25000# VSS 0.38174f $ **FLOATING
C1236 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.D VSS 0.4595f $ **FLOATING
C1237 a_61707_25000# VSS 0.36409f $ **FLOATING
C1238 3bit_freq_divider_1.freq_div_cell_0.Cin VSS 1.81006f $ **FLOATING
C1239 a_60967_24990# VSS 0.27856f $ **FLOATING
C1240 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.Q VSS 2.27033f $ **FLOATING
C1241 a_60584_24580# VSS 0.16608f $ **FLOATING
C1242 a_60385_24947# VSS 0.21087f $ **FLOATING
C1243 a_56137_24678# VSS 0.21087f $ **FLOATING
C1244 3bit_freq_divider_1.sg13g2_tiehi_1.L_HI VSS 1.60229f $ **FLOATING
C1245 a_60385_24717# VSS 0.17977f $ **FLOATING
C1246 a_60479_25023# VSS 0.01118f $ **FLOATING
C1247 a_55941_24882# VSS 0.16608f $ **FLOATING
C1248 3bit_freq_divider_0.dff_nclk_0.nRST VSS 1.20799f $ **FLOATING
C1249 a_51622_24863# VSS 0.17085f $ **FLOATING
C1250 3bit_freq_divider_0.freq_div_cell_0.Cin VSS 1.81006f $ **FLOATING
C1251 a_55345_24897# VSS 0.27856f $ **FLOATING
C1252 a_56039_25022# VSS 0.01118f $ **FLOATING
C1253 a_56013_24979# VSS 0.17977f $ **FLOATING
C1254 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.D VSS 0.4595f $ **FLOATING
C1255 a_54434_24904# VSS 0.36409f $ **FLOATING
C1256 3bit_freq_divider_0.sg13g2_or3_1_0.C VSS 2.00844f $ **FLOATING
C1257 a_52065_24890# VSS 0.01158f $ **FLOATING
C1258 a_51721_24988# VSS 0.21807f $ **FLOATING
C1259 a_51759_25014# VSS 0.18902f $ **FLOATING
C1260 a_52886_24904# VSS 0.38144f $ **FLOATING
C1261 3bit_freq_divider_0.sg13g2_tiehi_1.L_HI VSS 1.60229f $ **FLOATING
C1262 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.Q VSS 2.27033f $ **FLOATING
C1263 a_47954_28913# VSS 0.97627f $ **FLOATING
C1264 a_46817_27899# VSS 1.26528f $ **FLOATING
C1265 a_45658_27900# VSS 1.24513f $ **FLOATING
C1266 PFD_0.VCO_CLK VSS 5.09845f $ **FLOATING
C1267 a_48909_28913# VSS 1.03223f $ **FLOATING
C1268 a_45451_28860# VSS 1.00878f $ **FLOATING
C1269 a_47777_29803# VSS 1.2524f $ **FLOATING
C1270 a_46749_30782# VSS 1.31435f $ **FLOATING
C1271 a_45579_29803# VSS 0.97532f $ **FLOATING
C1272 a_59799_40285# VSS 0.05072f $ **FLOATING
C1273 a_58453_40283# VSS 0.04654f $ **FLOATING
C1274 a_57111_40283# VSS 0.0474f $ **FLOATING
C1275 a_55769_40283# VSS 0.04814f $ **FLOATING
C1276 a_54427_40283# VSS 0.04567f $ **FLOATING
C1277 a_53085_40283# VSS 0.07408f $ **FLOATING
C1278 a_58515_40413# VSS 4.51596f $ **FLOATING
C1279 a_57173_40413# VSS 4.66235f $ **FLOATING
C1280 a_55831_40413# VSS 4.71205f $ **FLOATING
C1281 a_54489_40413# VSS 5.15226f $ **FLOATING
C1282 a_53147_40413# VSS 5.26745f $ **FLOATING
C1283 a_59800_40852# VSS 0.75306f $ **FLOATING
C1284 a_58454_40850# VSS 0.8045f $ **FLOATING
C1285 a_57112_40850# VSS 0.81785f $ **FLOATING
C1286 a_55770_40850# VSS 0.82955f $ **FLOATING
C1287 a_54428_40850# VSS 0.82862f $ **FLOATING
C1288 a_53086_40850# VSS 0.83893f $ **FLOATING
C1289 a_58653_42591# VSS 0.65187f $ **FLOATING
C1290 a_57311_42591# VSS 0.67139f $ **FLOATING
C1291 a_55969_42591# VSS 0.6715f $ **FLOATING
C1292 a_54627_42591# VSS 0.67644f $ **FLOATING
C1293 a_53285_42591# VSS 0.68389f $ **FLOATING
C1294 3bit_freq_divider_0.CLK_IN VSS 20.6212f $ **FLOATING
C1295 a_57178_43159# VSS 5.00808f $ **FLOATING
C1296 a_55836_43159# VSS 4.39926f $ **FLOATING
C1297 a_54494_43159# VSS 4.398f $ **FLOATING
C1298 a_53152_43159# VSS 4.66518f $ **FLOATING
C1299 a_52944_43077# VSS 6.1695f $ **FLOATING
C1300 a_58426_43159# VSS 0.05888f $ **FLOATING
C1301 a_57084_43159# VSS 0.03844f $ **FLOATING
C1302 a_55742_43159# VSS 0.04051f $ **FLOATING
C1303 a_54400_43159# VSS 0.04084f $ **FLOATING
C1304 a_53058_43159# VSS 0.05472f $ **FLOATING
C1305 a_53022_43738# VSS 5.68098f $ **FLOATING
C1306 a_54747_49259# VSS 0.16684f $ **FLOATING
C1307 PFD_0.DOWN VSS 13.9137f $ **FLOATING
C1308 a_60528_49446# VSS 0.16044f
C1309 a_56695_49467# VSS 0.14015f
C1310 vco_wob_0.vctl VSS 17.2852f $ **FLOATING
C1311 a_56887_49467# VSS 8.04158f $ **FLOATING
C1312 a_54357_49278# VSS 0.26592f $ **FLOATING
C1313 PFD_0.UP VSS 12.6721f $ **FLOATING
C1314 charge_pump_0.vout VSS 28.7608f $ **FLOATING
C1315 a_56828_53480# VSS 2.32258f
C1316 a_56742_53480# VSS 1.67237f $ **FLOATING
C1317 a_59097_54704# VSS 0.1681f $ **FLOATING
C1318 a_58536_54976# VSS 0.61525f $ **FLOATING
C1319 a_58734_56203# VSS 0.05948f $ **FLOATING
C1320 charge_pump_0.bias_p VSS 5.47872f $ **FLOATING
C1321 charge_pump_0.bias_n VSS 6.55127f $ **FLOATING
C1322 3bit_freq_divider_0.EN VSS 51.6717f $ **FLOATING
C1323 a_55948_56737# VSS 1.95792f
C1324 a_55862_56737# VSS 0.99714f $ **FLOATING
.ends
