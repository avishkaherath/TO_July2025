* Extracted by KLayout with SG13G2 LVS runset on : 02/09/2025 10:55

.SUBCKT FMD_QNC_PLL_3BIT_DIV
X$1 \$1 \$1 \$44 \$2 \$39 \$42 \$11 \$11 Bias_gen
X$29517 \$1 \$11 \$12 \$13 \$41 \$15 PFD
X$37272 \$11 \$1 \$44 \$2 sg13g2_inv_1
X$38503 \$1 \$40 \$30 loop_filter
X$42292 \$I90878 \$11 \$1 sg13g2_tiehi
X$42293 \$I90873 \$I90877 \$I90877 \$13 \$1 \$I90878 \$11 dff_nclk
X$42294 \$11 \$1 \$I90875 \$I90876 \$I90874 \$I90873 sg13g2_or3_1
X$42295 \$I90880 \$I90879 \$I90872 \$7 \$I90874 \$1 \$I90873 \$11 freq_div_cell
X$42296 \$I90881 \$I90880 \$I90872 \$8 \$I90875 \$1 \$I90873 \$11 freq_div_cell
X$42297 \$I90881 \$11 \$1 sg13g2_tiehi
X$42298 \$I90879 \$I90882 \$I90872 \$6 \$I90876 \$1 \$I90873 \$11 freq_div_cell
X$42299 \$11 \$1 \$I90872 \$4 \$2 sg13g2_nand2_1
X$42300 \$I90889 \$11 \$1 sg13g2_tiehi
X$42301 \$I90884 \$I90888 \$I90888 \$10 \$1 \$I90889 \$11 dff_nclk
X$42302 \$11 \$1 \$I90886 \$I90887 \$I90885 \$I90884 sg13g2_or3_1
X$42303 \$I90891 \$I90890 \$I90883 \$9 \$I90885 \$1 \$I90884 \$11 freq_div_cell
X$42304 \$I90892 \$I90891 \$I90883 \$14 \$I90886 \$1 \$I90884 \$11 freq_div_cell
X$42305 \$I90892 \$11 \$1 sg13g2_tiehi
X$42306 \$I90890 \$I90893 \$I90883 \$5 \$I90887 \$1 \$I90884 \$11 freq_div_cell
X$42307 \$11 \$1 \$I90883 \$4 \$2 sg13g2_nand2_1
M$1 \$1 \$39 \$I42161 \$1 sg13_lv_nmos L=0.13u W=1.2u AS=0.408p AD=0.228p
+ PS=3.08u PD=1.58u
M$2 \$I42161 \$12 \$40 \$1 sg13_lv_nmos L=0.13u W=1.2u AS=0.228p AD=0.408p
+ PS=1.58u PD=3.08u
M$3 \$40 \$I42160 \$43 \$11 sg13_lv_pmos L=0.13u W=0.15u AS=0.1005p AD=0.0555p
+ PS=1.34u PD=0.74u
M$4 \$43 \$42 \$11 \$11 sg13_lv_pmos L=0.13u W=0.15u AS=0.0555p AD=0.1005p
+ PS=0.74u PD=1.34u
M$5 \$28 \$23 \$24 \$1 sg13_lv_nmos L=0.13u W=1u AS=0.28p AD=0.28p PS=2.62u
+ PD=2.62u
M$7 \$1 \$30 \$I90853 \$1 sg13_lv_nmos L=0.13u W=0.6u AS=0.159p AD=0.159p
+ PS=1.96u PD=1.96u
M$9 \$1 \$30 \$27 \$1 sg13_lv_nmos L=0.13u W=0.6u AS=0.159p AD=0.159p PS=1.96u
+ PD=1.96u
M$11 \$1 \$30 \$I90855 \$1 sg13_lv_nmos L=0.13u W=0.6u AS=0.159p AD=0.159p
+ PS=1.96u PD=1.96u
M$13 \$1 \$30 \$I90856 \$1 sg13_lv_nmos L=0.13u W=0.6u AS=0.159p AD=0.159p
+ PS=1.96u PD=1.96u
M$15 \$27 \$25 \$26 \$1 sg13_lv_nmos L=0.13u W=1u AS=0.28p AD=0.28p PS=2.62u
+ PD=2.62u
M$17 \$1 \$30 \$I90857 \$1 sg13_lv_nmos L=0.13u W=0.6u AS=0.159p AD=0.159p
+ PS=1.96u PD=1.96u
M$19 \$I90852 \$22 \$23 \$1 sg13_lv_nmos L=0.13u W=1u AS=0.28p AD=0.28p
+ PS=2.62u PD=2.62u
M$21 \$I90851 \$24 \$25 \$1 sg13_lv_nmos L=0.13u W=1u AS=0.28p AD=0.28p
+ PS=2.62u PD=2.62u
M$23 \$I90853 \$4 \$22 \$1 sg13_lv_nmos L=0.13u W=1u AS=0.265p AD=0.265p
+ PS=2.56u PD=2.56u
M$25 \$1 \$30 \$I90851 \$1 sg13_lv_nmos L=0.13u W=0.6u AS=0.159p AD=0.159p
+ PS=1.96u PD=1.96u
M$27 \$1 \$30 \$28 \$1 sg13_lv_nmos L=0.13u W=0.6u AS=0.159p AD=0.159p PS=1.96u
+ PD=1.96u
M$29 \$1 \$30 \$I90858 \$1 sg13_lv_nmos L=0.13u W=0.6u AS=0.159p AD=0.159p
+ PS=1.96u PD=1.96u
M$31 \$1 \$30 \$I90854 \$1 sg13_lv_nmos L=0.13u W=0.6u AS=0.159p AD=0.159p
+ PS=1.96u PD=1.96u
M$33 \$1 \$30 \$16 \$1 sg13_lv_nmos L=0.13u W=0.6u AS=0.159p AD=0.159p PS=1.96u
+ PD=1.96u
M$35 \$1 \$30 \$I90850 \$1 sg13_lv_nmos L=0.13u W=0.6u AS=0.159p AD=0.159p
+ PS=1.96u PD=1.96u
M$37 \$1 \$30 \$I90852 \$1 sg13_lv_nmos L=0.13u W=0.6u AS=0.159p AD=0.159p
+ PS=1.96u PD=1.96u
M$39 \$I90850 \$26 \$I90849 \$1 sg13_lv_nmos L=0.13u W=1u AS=0.28p AD=0.28p
+ PS=2.62u PD=2.62u
M$41 \$11 \$16 \$I90843 \$11 sg13_lv_pmos L=0.13u W=0.8u AS=0.28325p
+ AD=0.28175p PS=3.575u PD=3.565u
M$45 \$I90846 \$4 \$22 \$11 sg13_lv_pmos L=0.13u W=2u AS=0.455p AD=0.455p
+ PS=4.32u PD=4.32u
M$49 \$11 \$16 \$16 \$11 sg13_lv_pmos L=0.13u W=0.8u AS=0.2825p AD=0.2825p
+ PS=3.57u PD=3.57u
M$53 \$11 \$16 \$I90864 \$11 sg13_lv_pmos L=0.13u W=0.8u AS=0.23825p
+ AD=0.32675p PS=2.975u PD=4.165u
M$57 \$11 \$16 \$I90847 \$11 sg13_lv_pmos L=0.13u W=0.8u AS=0.28325p
+ AD=0.28175p PS=3.575u PD=3.565u
M$61 \$11 \$16 \$I90863 \$11 sg13_lv_pmos L=0.13u W=0.8u AS=0.23825p
+ AD=0.32675p PS=2.975u PD=4.165u
M$65 \$I90845 \$22 \$23 \$11 sg13_lv_pmos L=0.13u W=2u AS=0.455p AD=0.455p
+ PS=4.32u PD=4.32u
M$69 \$I90847 \$26 \$I90849 \$11 sg13_lv_pmos L=0.13u W=2u AS=0.455p AD=0.455p
+ PS=4.32u PD=4.32u
M$73 \$11 \$16 \$I90844 \$11 sg13_lv_pmos L=0.13u W=0.8u AS=0.28325p
+ AD=0.28175p PS=3.575u PD=3.565u
M$77 \$I90843 \$24 \$25 \$11 sg13_lv_pmos L=0.13u W=2u AS=0.455p AD=0.455p
+ PS=4.32u PD=4.32u
M$81 \$I90848 \$25 \$26 \$11 sg13_lv_pmos L=0.13u W=2u AS=0.455p AD=0.455p
+ PS=4.32u PD=4.32u
M$85 \$11 \$16 \$I90845 \$11 sg13_lv_pmos L=0.13u W=0.8u AS=0.28325p
+ AD=0.28175p PS=3.575u PD=3.565u
M$89 \$11 \$16 \$I90846 \$11 sg13_lv_pmos L=0.13u W=0.8u AS=0.281p AD=0.281p
+ PS=3.56u PD=3.56u
M$93 \$11 \$16 \$I90848 \$11 sg13_lv_pmos L=0.13u W=0.8u AS=0.28325p
+ AD=0.28175p PS=3.575u PD=3.565u
M$97 \$11 \$16 \$I90865 \$11 sg13_lv_pmos L=0.13u W=0.8u AS=0.23825p
+ AD=0.32675p PS=2.975u PD=4.165u
M$101 \$11 \$16 \$I90862 \$11 sg13_lv_pmos L=0.13u W=0.8u AS=0.23825p
+ AD=0.32675p PS=2.975u PD=4.165u
M$105 \$11 \$16 \$I90866 \$11 sg13_lv_pmos L=0.13u W=0.8u AS=0.23825p
+ AD=0.32675p PS=2.975u PD=4.165u
M$109 \$I90844 \$23 \$24 \$11 sg13_lv_pmos L=0.13u W=2u AS=0.455p AD=0.455p
+ PS=4.32u PD=4.32u
M$113 \$I42160 \$41 \$11 \$11 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.102p
+ PS=1.28u PD=1.28u
M$114 \$1 \$41 \$I42160 \$1 sg13_lv_nmos L=0.13u W=0.15u AS=0.1005p AD=0.1005p
+ PS=1.34u PD=1.34u
C$115 \$25 \$1 cap_cmim w=6.99u l=6.99u A=48.8601p P=27.96u m=1
C$116 \$24 \$1 cap_cmim w=6.99u l=6.99u A=48.8601p P=27.96u m=1
C$117 \$33 \$1 cap_cmim w=6.99u l=6.99u A=48.8601p P=27.96u m=1
C$118 \$I90859 \$1 cap_cmim w=6.99u l=6.99u A=48.8601p P=27.96u m=1
C$119 \$I90849 \$1 cap_cmim w=6.99u l=6.99u A=48.8601p P=27.96u m=1
C$120 \$26 \$1 cap_cmim w=6.99u l=6.99u A=48.8601p P=27.96u m=1
C$121 \$23 \$1 cap_cmim w=6.99u l=6.99u A=48.8601p P=27.96u m=1
C$122 \$22 \$1 cap_cmim w=6.99u l=6.99u A=48.8601p P=27.96u m=1
C$123 \$I90861 \$1 cap_cmim w=6.99u l=6.99u A=48.8601p P=27.96u m=1
C$124 \$4 \$1 cap_cmim w=6.99u l=6.99u A=48.8601p P=27.96u m=1
C$125 \$I90860 \$1 cap_cmim w=6.99u l=6.99u A=48.8601p P=27.96u m=1
M$126 \$I90854 \$I90849 \$33 \$1 sg13_lv_nmos L=0.13u W=1u AS=0.265p AD=0.265p
+ PS=2.56u PD=2.56u
M$128 \$I90862 \$I90849 \$33 \$11 sg13_lv_pmos L=0.13u W=2u AS=0.455p AD=0.455p
+ PS=4.32u PD=4.32u
M$132 \$I90855 \$33 \$I90868 \$1 sg13_lv_nmos L=0.13u W=1u AS=0.265p AD=0.265p
+ PS=2.56u PD=2.56u
M$134 \$I90863 \$33 \$I90859 \$11 sg13_lv_pmos L=0.13u W=2u AS=0.455p AD=0.455p
+ PS=4.32u PD=4.32u
M$138 \$I90857 \$I90859 \$I90870 \$1 sg13_lv_nmos L=0.13u W=1u AS=0.265p
+ AD=0.265p PS=2.56u PD=2.56u
M$140 \$I90864 \$I90859 \$I90860 \$11 sg13_lv_pmos L=0.13u W=2u AS=0.455p
+ AD=0.455p PS=4.32u PD=4.32u
M$144 \$I90858 \$I90860 \$I90871 \$1 sg13_lv_nmos L=0.13u W=1u AS=0.265p
+ AD=0.265p PS=2.56u PD=2.56u
M$146 \$I90865 \$I90860 \$I90861 \$11 sg13_lv_pmos L=0.13u W=2u AS=0.455p
+ AD=0.455p PS=4.32u PD=4.32u
M$150 \$I90856 \$I90861 \$I90869 \$1 sg13_lv_nmos L=0.13u W=1u AS=0.265p
+ AD=0.265p PS=2.56u PD=2.56u
M$152 \$I90866 \$I90861 \$4 \$11 sg13_lv_pmos L=0.13u W=2u AS=0.455p AD=0.455p
+ PS=4.32u PD=4.32u
.ENDS FMD_QNC_PLL_3BIT_DIV

.SUBCKT PFD VSS VDD DOWN VCO_CLK UP Ref_CLK
M$1 \$5 VCO_CLK \$7 VSS sg13_lv_nmos L=0.15u W=0.84u AS=0.2226p AD=0.2226p
+ PS=2.32u PD=2.32u
M$3 \$10 Ref_CLK \$12 VSS sg13_lv_nmos L=0.15u W=0.84u AS=0.2226p AD=0.2226p
+ PS=2.32u PD=2.32u
M$5 VSS \$13 UP VSS sg13_lv_nmos L=0.15u W=0.48u AS=0.1632p AD=0.1632p PS=1.64u
+ PD=1.64u
M$6 VSS \$4 DOWN VSS sg13_lv_nmos L=0.15u W=0.48u AS=0.1632p AD=0.1632p
+ PS=1.64u PD=1.64u
M$7 \$8 VCO_CLK VSS VSS sg13_lv_nmos L=0.15u W=0.36u AS=0.1224p AD=0.1224p
+ PS=1.4u PD=1.4u
M$8 VSS \$10 \$13 VSS sg13_lv_nmos L=0.15u W=0.36u AS=0.1224p AD=0.1224p
+ PS=1.4u PD=1.4u
M$9 VSS \$5 \$4 VSS sg13_lv_nmos L=0.15u W=0.36u AS=0.1224p AD=0.1224p PS=1.4u
+ PD=1.4u
M$10 \$9 Ref_CLK VSS VSS sg13_lv_nmos L=0.15u W=0.36u AS=0.1224p AD=0.1224p
+ PS=1.4u PD=1.4u
M$11 VDD \$13 UP VDD sg13_lv_pmos L=0.15u W=0.96u AS=0.2304p AD=0.2304p
+ PS=2.72u PD=2.72u
M$14 VDD \$4 DOWN VDD sg13_lv_pmos L=0.15u W=0.96u AS=0.2304p AD=0.2304p
+ PS=2.72u PD=2.72u
M$17 \$13 \$10 VDD VDD sg13_lv_pmos L=0.15u W=0.72u AS=0.1908p AD=0.1908p
+ PS=2.14u PD=2.14u
M$19 VDD \$5 \$4 VDD sg13_lv_pmos L=0.15u W=0.72u AS=0.1908p AD=0.1908p
+ PS=2.14u PD=2.14u
M$21 \$8 Ref_CLK \$12 VSS sg13_lv_nmos L=0.15u W=1.8u AS=0.396p AD=0.396p
+ PS=4.36u PD=4.36u
M$26 \$9 VCO_CLK \$7 VSS sg13_lv_nmos L=0.15u W=1.8u AS=0.396p AD=0.396p
+ PS=4.36u PD=4.36u
M$31 \$12 Ref_CLK VDD VDD sg13_lv_pmos L=0.15u W=0.64u AS=0.1696p AD=0.1696p
+ PS=2.02u PD=2.02u
M$33 \$7 VCO_CLK VDD VDD sg13_lv_pmos L=0.15u W=0.64u AS=0.1696p AD=0.1696p
+ PS=2.02u PD=2.02u
M$35 \$5 VCO_CLK VCO_CLK VDD sg13_lv_pmos L=0.15u W=0.64u AS=0.1696p AD=0.1696p
+ PS=2.02u PD=2.02u
M$37 \$10 Ref_CLK Ref_CLK VDD sg13_lv_pmos L=0.15u W=0.64u AS=0.1696p
+ AD=0.1696p PS=2.02u PD=2.02u
.ENDS PFD

.SUBCKT Bias_gen \$1 \$2 enb en \$6 \$9 \$10 \$13
R$1 \$11 \$13 rhigh w=1u l=12u ps=0 b=0 m=1
R$2 \$3 \$2 rhigh w=1u l=12u ps=0 b=0 m=1
M$3 \$7 \$6 \$2 \$1 sg13_lv_nmos L=1u W=1u AS=0.34p AD=0.34p PS=2.68u PD=2.68u
M$4 \$9 \$6 \$3 \$1 sg13_lv_nmos L=1u W=1u AS=0.34p AD=0.34p PS=2.68u PD=2.68u
M$5 \$6 \$6 \$2 \$1 sg13_lv_nmos L=1u W=1u AS=0.34p AD=0.34p PS=2.68u PD=2.68u
M$6 \$9 \$7 \$8 \$1 sg13_lv_nmos L=0.15u W=0.5u AS=0.17p AD=0.17p PS=1.68u
+ PD=1.68u
M$7 \$6 enb \$2 \$1 sg13_lv_nmos L=0.15u W=0.5u AS=0.17p AD=0.17p PS=1.68u
+ PD=1.68u
M$8 \$8 en \$2 \$1 sg13_lv_nmos L=0.15u W=0.5u AS=0.17p AD=0.17p PS=1.68u
+ PD=1.68u
M$9 \$6 \$9 \$11 \$10 sg13_lv_pmos L=1u W=4u AS=1.06p AD=1.06p PS=7.06u PD=7.06u
M$11 \$13 \$9 \$9 \$10 sg13_lv_pmos L=1u W=2u AS=0.68p AD=0.68p PS=4.68u
+ PD=4.68u
M$12 \$13 \$12 \$12 \$10 sg13_lv_pmos L=0.15u W=0.5u AS=0.17p AD=0.17p PS=1.68u
+ PD=1.68u
M$13 \$13 en \$9 \$10 sg13_lv_pmos L=0.15u W=0.5u AS=0.17p AD=0.17p PS=1.68u
+ PD=1.68u
M$14 \$12 \$7 \$7 \$10 sg13_lv_pmos L=0.15u W=0.5u AS=0.17p AD=0.17p PS=1.68u
+ PD=1.68u
M$15 \$13 en \$7 \$10 sg13_lv_pmos L=0.15u W=0.5u AS=0.17p AD=0.17p PS=1.68u
+ PD=1.68u
.ENDS Bias_gen

.SUBCKT loop_filter \$1 \$2 \$3
M$1 \$1 \$2 \$1 \$1 sg13_lv_nmos L=0.65u W=45u AS=9p AD=9p PS=60u PD=60u
R$31 \$2 \$3 rhigh w=0.6u l=0.96u ps=0 b=0 m=1
R$32 \$4 \$2 rhigh w=0.5u l=0.96u ps=0 b=0 m=1
M$33 \$1 \$3 \$1 \$1 sg13_lv_nmos L=0.13u W=0.3u AS=0.201p AD=0.201p PS=2.68u
+ PD=2.68u
M$35 \$1 \$4 \$1 \$1 sg13_lv_nmos L=0.65u W=15u AS=3p AD=3p PS=28u PD=28u
.ENDS loop_filter

.SUBCKT sg13g2_nand2_1 VDD VSS Y A B
M$1 VSS B \$6 VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.2516p AD=0.0666p PS=2.16u
+ PD=0.92u
M$2 \$6 A Y VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.0666p AD=0.2516p PS=0.92u
+ PD=2.16u
M$3 VDD B Y VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.3808p AD=0.2128p PS=2.92u
+ PD=1.5u
M$4 Y A VDD VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.2128p AD=0.3808p PS=1.5u
+ PD=2.92u
.ENDS sg13g2_nand2_1

.SUBCKT sg13g2_or3_1 VDD VSS C A B X
M$1 \$6 C VSS VSS sg13_lv_nmos L=0.13u W=0.55u AS=0.187p AD=0.1045p PS=1.78u
+ PD=0.93u
M$2 VSS B \$6 VSS sg13_lv_nmos L=0.13u W=0.55u AS=0.1045p AD=0.198p PS=0.93u
+ PD=1.27u
M$3 \$6 A VSS VSS sg13_lv_nmos L=0.13u W=0.55u AS=0.198p AD=0.13395p PS=1.27u
+ PD=1.12u
M$4 VSS \$6 X VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.13395p AD=0.2516p PS=1.12u
+ PD=2.16u
M$5 \$6 C \$9 VDD sg13_lv_pmos L=0.13u W=1u AS=0.34p AD=0.1275p PS=2.68u
+ PD=1.255u
M$6 \$9 B \$8 VDD sg13_lv_pmos L=0.13u W=1u AS=0.1275p AD=0.22p PS=1.255u
+ PD=1.44u
M$7 \$8 A VDD VDD sg13_lv_pmos L=0.13u W=1u AS=0.22p AD=0.3822p PS=1.44u
+ PD=1.84u
M$8 VDD \$6 X VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.3822p AD=0.3808p PS=1.84u
+ PD=2.92u
.ENDS sg13g2_or3_1

.SUBCKT sg13g2_tiehi L_HI VDD VSS
M$1 VSS \$4 \$4 VSS sg13_lv_nmos L=0.13u W=0.3u AS=0.2307p AD=0.102p PS=1.615u
+ PD=1.28u
M$2 VSS \$3 \$1 VSS sg13_lv_nmos L=0.13u W=0.795u AS=0.2307p AD=0.274275p
+ PS=1.615u PD=2.28u
M$3 \$3 \$4 VDD VDD sg13_lv_pmos L=0.13u W=0.66u AS=0.2442p AD=0.4657125p
+ PS=2.06u PD=2.54u
M$4 VDD \$1 L_HI VDD sg13_lv_pmos L=0.13u W=1.155u AS=0.4657125p AD=0.3927p
+ PS=2.54u PD=2.99u
.ENDS sg13g2_tiehi

.SUBCKT freq_div_cell Cin Cout CLK BIT DIV \$7 nRST \$11
X$1 Cin \$6 \$9 Cout \$7 \$11 half_add
X$2 CLK \$9 \$I8 \$6 \$7 nRST \$11 dff_nclk
X$3 \$7 DIV \$11 \$6 BIT sg13g2_xor2_1
.ENDS freq_div_cell

.SUBCKT dff_nclk nCLK D nQ Q \$6 nRST \$9
X$1 \$9 \$6 nCLK \$5 sg13g2_inv_1
X$2 \$6 nRST nQ Q D \$5 \$9 sg13g2_dfrbp_1
.ENDS dff_nclk

.SUBCKT half_add inA inB sum cout \$5 \$6
X$1 \$5 sum \$6 inA inB sg13g2_xor2_1
X$2 \$6 \$5 cout inA inB sg13g2_and2_1
.ENDS half_add

.SUBCKT sg13g2_dfrbp_1 VSS RESET_B Q_N Q D CLK VDD
M$1 \$5 \$11 \$19 VSS sg13_lv_nmos L=0.13u W=0.42u AS=0.2017p AD=0.0546p
+ PS=1.48u PD=0.68u
M$2 \$19 \$6 VSS VSS sg13_lv_nmos L=0.13u W=0.42u AS=0.0546p AD=0.0903p
+ PS=0.68u PD=0.85u
M$3 VSS RESET_B \$18 VSS sg13_lv_nmos L=0.13u W=0.42u AS=0.0903p AD=0.04725p
+ PS=0.85u PD=0.645u
M$4 \$18 \$5 \$6 VSS sg13_lv_nmos L=0.13u W=0.42u AS=0.04725p AD=0.1428p
+ PS=0.645u PD=1.52u
M$5 VSS \$13 \$14 VSS sg13_lv_nmos L=0.13u W=0.64u AS=0.1825p AD=0.193975p
+ PS=1.325u PD=1.29u
M$6 \$14 \$3 \$5 VSS sg13_lv_nmos L=0.13u W=0.64u AS=0.193975p AD=0.2017p
+ PS=1.29u PD=1.48u
M$7 \$4 \$11 \$13 VSS sg13_lv_nmos L=0.13u W=0.42u AS=0.1428p AD=0.0798p
+ PS=1.52u PD=0.8u
M$8 \$13 \$3 \$16 VSS sg13_lv_nmos L=0.13u W=0.42u AS=0.0798p AD=0.0546p
+ PS=0.8u PD=0.68u
M$9 \$16 \$14 \$17 VSS sg13_lv_nmos L=0.13u W=0.42u AS=0.0546p AD=0.0483p
+ PS=0.68u PD=0.65u
M$10 VSS RESET_B \$17 VSS sg13_lv_nmos L=0.13u W=0.42u AS=0.1825p AD=0.0483p
+ PS=1.325u PD=0.65u
M$11 \$8 \$5 VSS VSS sg13_lv_nmos L=0.13u W=0.55u AS=0.187p AD=0.14505p
+ PS=1.78u PD=1.15u
M$12 VSS \$8 Q VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.14505p AD=0.2516p PS=1.15u
+ PD=2.16u
M$13 VSS \$5 Q_N VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.2516p AD=0.2775p
+ PS=2.16u PD=2.23u
M$14 VSS CLK \$11 VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.1544p AD=0.2516p
+ PS=1.235u PD=2.16u
M$15 VSS \$11 \$3 VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.1544p AD=0.2516p
+ PS=1.235u PD=2.16u
M$16 \$4 D \$15 VSS sg13_lv_nmos L=0.13u W=0.42u AS=0.1428p AD=0.0504p PS=1.52u
+ PD=0.66u
M$17 \$15 RESET_B VSS VSS sg13_lv_nmos L=0.13u W=0.42u AS=0.0504p AD=0.1428p
+ PS=0.66u PD=1.52u
M$18 VDD \$13 \$14 VDD sg13_lv_pmos L=0.13u W=1u AS=0.34p AD=0.19p PS=2.68u
+ PD=1.38u
M$19 \$14 \$11 \$5 VDD sg13_lv_pmos L=0.13u W=1u AS=0.19p AD=0.17695p PS=1.38u
+ PD=1.56u
M$20 \$5 \$3 \$22 VDD sg13_lv_pmos L=0.13u W=0.42u AS=0.17695p AD=0.04305p
+ PS=1.56u PD=0.625u
M$21 \$22 \$6 VDD VDD sg13_lv_pmos L=0.13u W=0.42u AS=0.04305p AD=0.0798p
+ PS=0.625u PD=0.8u
M$22 VDD RESET_B \$6 VDD sg13_lv_pmos L=0.13u W=0.42u AS=0.0798p AD=0.0798p
+ PS=0.8u PD=0.8u
M$23 VDD \$5 \$6 VDD sg13_lv_pmos L=0.13u W=0.42u AS=0.2163p AD=0.0798p
+ PS=1.55u PD=0.8u
M$24 VDD \$5 Q_N VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.2163p AD=0.7616p
+ PS=1.55u PD=3.6u
M$25 \$4 \$3 \$13 VDD sg13_lv_pmos L=0.13u W=0.42u AS=0.1428p AD=0.0798p
+ PS=1.52u PD=0.8u
M$26 \$13 \$11 \$21 VDD sg13_lv_pmos L=0.13u W=0.42u AS=0.0798p AD=0.05145p
+ PS=0.8u PD=0.665u
M$27 \$21 \$14 VDD VDD sg13_lv_pmos L=0.13u W=0.42u AS=0.05145p AD=0.11785p
+ PS=0.665u PD=1.025u
M$28 VDD RESET_B \$13 VDD sg13_lv_pmos L=0.13u W=0.42u AS=0.11785p AD=0.1533p
+ PS=1.025u PD=1.57u
M$29 \$11 CLK VDD VDD sg13_lv_pmos L=0.13u W=1u AS=0.34p AD=0.19p PS=2.68u
+ PD=1.38u
M$30 VDD \$11 \$3 VDD sg13_lv_pmos L=0.13u W=1u AS=0.19p AD=0.34p PS=1.38u
+ PD=2.68u
M$31 VDD D \$4 VDD sg13_lv_pmos L=0.13u W=0.42u AS=0.1428p AD=0.0798p PS=1.52u
+ PD=0.8u
M$32 \$4 RESET_B VDD VDD sg13_lv_pmos L=0.13u W=0.42u AS=0.0798p AD=0.1428p
+ PS=0.8u PD=1.52u
M$33 VDD \$5 \$8 VDD sg13_lv_pmos L=0.13u W=0.84u AS=0.2016p AD=0.2856p PS=1.5u
+ PD=2.36u
M$34 VDD \$8 Q VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.2016p AD=0.3808p PS=1.5u
+ PD=2.92u
.ENDS sg13g2_dfrbp_1

.SUBCKT sg13g2_inv_1 VDD VSS A Y
M$1 VSS A Y VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.259p AD=0.259p PS=2.18u
+ PD=2.18u
M$2 VDD A Y VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.392p AD=0.392p PS=2.94u
+ PD=2.94u
.ENDS sg13g2_inv_1

.SUBCKT sg13g2_and2_1 VDD VSS X A B
M$1 \$6 A \$7 VSS sg13_lv_nmos L=0.13u W=0.64u AS=0.2176p AD=0.1216p PS=1.96u
+ PD=1.02u
M$2 VSS B \$7 VSS sg13_lv_nmos L=0.13u W=0.64u AS=0.1331p AD=0.1216p PS=1.12u
+ PD=1.02u
M$3 VSS \$6 X VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.1331p AD=0.2516p PS=1.12u
+ PD=2.16u
M$4 VDD A \$6 VDD sg13_lv_pmos L=0.13u W=0.84u AS=0.2856p AD=0.1596p PS=2.36u
+ PD=1.22u
M$5 VDD B \$6 VDD sg13_lv_pmos L=0.13u W=0.84u AS=0.1918p AD=0.1596p PS=1.5u
+ PD=1.22u
M$6 VDD \$6 X VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.1918p AD=0.3808p PS=1.5u
+ PD=2.92u
.ENDS sg13g2_and2_1

.SUBCKT sg13g2_xor2_1 VSS X VDD A B
M$1 VSS A \$1 VSS sg13_lv_nmos L=0.13u W=0.55u AS=0.374p AD=0.174625p PS=2.46u
+ PD=1.185u
M$2 VSS B \$1 VSS sg13_lv_nmos L=0.13u W=0.55u AS=0.15245p AD=0.174625p
+ PS=1.17u PD=1.185u
M$3 VSS A \$8 VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.15245p AD=0.0888p PS=1.17u
+ PD=0.98u
M$4 \$8 B X VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.0888p AD=0.1628p PS=0.98u
+ PD=1.18u
M$5 X \$1 VSS VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.1628p AD=0.3108p PS=1.18u
+ PD=2.32u
M$6 \$3 A VDD VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.3808p AD=0.2128p PS=2.92u
+ PD=1.5u
M$7 VDD B \$3 VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.2128p AD=0.2128p PS=1.5u
+ PD=1.5u
M$8 \$3 \$1 X VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.2128p AD=0.3808p PS=1.5u
+ PD=2.92u
M$9 VDD A \$9 VDD sg13_lv_pmos L=0.13u W=1u AS=0.36p AD=0.1225p PS=2.72u
+ PD=1.245u
M$10 \$9 B \$1 VDD sg13_lv_pmos L=0.13u W=1u AS=0.1225p AD=0.34p PS=1.245u
+ PD=2.68u
.ENDS sg13g2_xor2_1
