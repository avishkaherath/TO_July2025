* NGSPICE file created from pll_3bitDiv.ext - technology: ihp-sg13g2

.subckt pll_3bitDiv CLK_IN CLK_OUT Y0 Y2 Y1 VDD VSS nEN X1 X2 X0
X0 VDD a_53968_20434# a_53899_20488# VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0.19p ps=1.38u w=1u l=0.13u
X1 VSS 3bit_freq_divider_1.dff_nclk_0.nCLK a_61488_20220# VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=50.4f ps=0.66u w=0.42u l=0.13u
X2 a_62119_20605# a_61691_20534# a_61394_20220# VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0.1428p ps=1.52u w=0.42u l=0.13u
X3 a_52924_22885# 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.Q VDD VDD sg13_lv_pmos ad=0.3808p pd=2.92u as=0.2128p ps=1.5u w=1.12u l=0.13u
X4 a_53065_20179# a_53738_20514# a_53702_20612# VDD sg13_lv_pmos ad=0.17695p pd=1.56u as=43.05f ps=0.625u w=0.42u l=0.13u
X5 a_62119_22361# 3bit_freq_divider_1.dff_nclk_0.nCLK VDD VDD sg13_lv_pmos ad=0.1533p pd=1.57u as=0.11785p ps=1.025u w=0.42u l=0.13u
X6 a_53152_43159# VSS cap_cmim l=6.99u w=6.99u
X7 VDD a_52950_22157# 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.Q VDD sg13_lv_pmos ad=0.2016p pd=1.5u as=0.3808p ps=2.92u w=1.12u l=0.13u
X8 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 3bit_freq_divider_1.sg13g2_nand2_1_0.Y VSS VSS sg13_lv_nmos ad=0.259p pd=2.18u as=0.259p ps=2.18u w=0.74u l=0.13u
X9 VSS 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.Q a_61061_23234# VSS sg13_lv_nmos ad=0.1331p pd=1.12u as=0.1216p ps=1.02u w=0.64u l=0.13u
X10 a_62879_24125# a_61887_24046# a_62654_23727# VDD sg13_lv_pmos ad=43.05f pd=0.625u as=0.17695p ps=1.56u w=0.42u l=0.13u
X11 a_53022_43738# a_53022_43738# VDD VDD sg13_lv_pmos ad=59f pd=0.74u as=0.104p ps=1.34u w=0.2u l=0.13u
X12 VSS a_55345_24897# 3bit_freq_divider_0.freq_div_cell_0.Cin VSS sg13_lv_nmos ad=0.1331p pd=1.12u as=0.2516p ps=2.16u w=0.74u l=0.13u
X13 a_64383_23434# a_64383_23628# VSS VSS sg13_lv_nmos ad=0.2516p pd=2.16u as=0.1544p ps=1.235u w=0.74u l=0.13u
X14 VDD a_53774_21934# a_53738_22270# VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0.34p ps=2.68u w=1u l=0.13u
X15 a_55485_23233# 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.Q VSS VSS sg13_lv_nmos ad=0.1216p pd=1.02u as=0.1331p ps=1.12u w=0.64u l=0.13u
X16 a_64383_23300# a_64383_23628# a_64424_22200# VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0.1428p ps=1.52u w=0.42u l=0.13u
X17 VSS charge_pump_0.vout VSS VSS sg13_lv_nmos ad=0.285p pd=1.88u as=0.53383n ps=1.58949m w=1.5u l=0.65u
X18 VDD a_53022_43738# a_57084_43159# VDD sg13_lv_pmos ad=0.104p pd=1.34u as=59f ps=0.74u w=0.2u l=0.13u
X19 VDD a_51648_21103# 3bit_freq_divider_0.dff_nclk_0.nCLK VDD sg13_lv_pmos ad=0.3822p pd=1.84u as=0.3808p ps=2.92u w=1.12u l=0.13u
X20 a_64383_23434# a_64383_23628# VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0.19p ps=1.38u w=1u l=0.13u
X21 a_54627_42591# vco_wob_0.vctl VSS VSS sg13_lv_nmos ad=65.99999f pd=0.74u as=0.102p ps=1.28u w=0.3u l=0.13u
X22 a_59799_40285# 3bit_freq_divider_0.CLK_IN a_58515_40413# VDD sg13_lv_pmos ad=0.17p pd=1.68u as=0.1106p ps=0.945u w=0.5u l=0.13u
X23 a_61972_23244# 3bit_freq_divider_1.freq_div_cell_0.Cin VSS VSS sg13_lv_nmos ad=88.8f pd=0.98u as=0.15245p ps=1.17u w=0.74u l=0.13u
X24 a_54494_43159# a_53152_43159# a_54627_42591# VSS sg13_lv_nmos ad=0.11p pd=0.94u as=0.17p ps=1.68u w=0.5u l=0.13u
X25 a_54427_40283# a_54489_40413# a_53147_40413# VDD sg13_lv_pmos ad=0.11p pd=0.94u as=0.11p ps=0.94u w=0.5u l=0.13u
X26 VDD 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.D a_54504_23771# VDD sg13_lv_pmos ad=0.1428p pd=1.52u as=79.8f ps=0.8u w=0.42u l=0.13u
X27 a_53774_20178# 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.sg13g2_dfrbp_1_0.CLK VSS VSS sg13_lv_nmos ad=0.2516p pd=2.16u as=0.1544p ps=1.235u w=0.74u l=0.13u
X28 a_54504_20259# 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.D a_55086_20219# VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=50.4f ps=0.66u w=0.42u l=0.13u
X29 charge_pump_0.bias_n charge_pump_0.bias_n VSS VSS sg13_lv_nmos ad=0.34p pd=2.68u as=0.34p ps=2.68u w=1u l=1u
X30 VSS 3bit_freq_divider_0.freq_div_cell_0.Cout a_54434_21392# VSS sg13_lv_nmos ad=0.374p pd=2.46u as=0.17462p ps=1.185u w=0.55u l=0.13u
X31 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.Q a_63463_23728# VSS VSS sg13_lv_nmos ad=0.2516p pd=2.16u as=0.14505p ps=1.15u w=0.74u l=0.13u
X32 a_47954_28913# PFD_0.VCO_CLK a_48909_28913# VSS sg13_lv_nmos ad=68.39999f pd=0.74u as=68.39999f ps=0.74u w=0.36u l=0.15u
X33 a_54898_21129# 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.Q a_54434_21392# VDD sg13_lv_pmos ad=0.1225p pd=1.245u as=0.34p ps=2.68u w=1u l=0.13u
X34 VSS charge_pump_0.vout VSS VSS sg13_lv_nmos ad=0.285p pd=1.88u as=0 ps=0 w=1.5u l=0.65u
X35 a_51693_23426# 3bit_freq_divider_0.dff_nclk_0.nRST VDD VDD sg13_lv_pmos ad=0.1533p pd=1.57u as=0.11785p ps=1.025u w=0.42u l=0.13u
X36 3bit_freq_divider_1.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 3bit_freq_divider_1.dff_nclk_0.nCLK VSS VSS sg13_lv_nmos ad=0.259p pd=2.18u as=0.259p ps=2.18u w=0.74u l=0.13u
X37 PFD_0.UP a_47777_29803# VSS VSS sg13_lv_nmos ad=0.1632p pd=1.64u as=0.1632p ps=1.64u w=0.48u l=0.15u
X38 VDD a_62654_23727# a_62900_23691# VDD sg13_lv_pmos ad=0.2163p pd=1.55u as=79.8f ps=0.8u w=0.42u l=0.13u
X39 a_54504_23771# 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.D a_55086_23731# VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=50.4f ps=0.66u w=0.42u l=0.13u
X40 a_60967_23234# 3bit_freq_divider_1.freq_div_cell_0.Cin VDD VDD sg13_lv_pmos ad=0.1596p pd=1.22u as=0.2856p ps=2.36u w=0.84u l=0.13u
X41 a_54602_23243# 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.Q 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.D VSS sg13_lv_nmos ad=88.8f pd=0.98u as=0.1628p ps=1.18u w=0.74u l=0.13u
X42 a_54898_24641# 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.Q a_54434_24904# VDD sg13_lv_pmos ad=0.1225p pd=1.245u as=0.34p ps=2.68u w=1u l=0.13u
X43 VDD 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.Q a_60967_21478# VDD sg13_lv_pmos ad=0.1918p pd=1.5u as=0.1596p ps=1.22u w=0.84u l=0.13u
X44 a_62221_24117# a_61691_24046# a_62119_24117# VDD sg13_lv_pmos ad=51.45f pd=0.665u as=79.8f ps=0.8u w=0.42u l=0.13u
X45 a_58426_43159# a_57178_43159# 3bit_freq_divider_0.CLK_IN VDD sg13_lv_pmos ad=0.11p pd=0.94u as=0.1106p ps=0.945u w=0.5u l=0.13u
X46 a_62246_20260# a_61887_20534# a_62119_20605# VSS sg13_lv_nmos ad=54.6f pd=0.68u as=79.8f ps=0.8u w=0.42u l=0.13u
X47 a_52074_23051# a_51684_22692# a_51693_23426# VSS sg13_lv_nmos ad=54.6f pd=0.68u as=79.8f ps=0.8u w=0.42u l=0.13u
X48 a_54504_22015# 3bit_freq_divider_0.dff_nclk_0.nCLK VDD VDD sg13_lv_pmos ad=79.8f pd=0.8u as=0.1428p ps=1.52u w=0.42u l=0.13u
X49 VDD a_55345_23141# 3bit_freq_divider_0.freq_div_cell_0.Cout VDD sg13_lv_pmos ad=0.1918p pd=1.5u as=0.3808p ps=2.92u w=1.12u l=0.13u
X50 a_64464_23130# a_64419_23326# a_64464_23052# VSS sg13_lv_nmos ad=48.3f pd=0.65u as=54.6f ps=0.68u w=0.42u l=0.13u
X51 VSS a_63255_21488# 3bit_freq_divider_1.sg13g2_or3_1_0.A VSS sg13_lv_nmos ad=0.3108p pd=2.32u as=0.1628p ps=1.18u w=0.74u l=0.13u
X52 a_61675_22886# 3bit_freq_divider_1.freq_div_cell_0.Cin VDD VDD sg13_lv_pmos ad=0.1225p pd=1.245u as=0.36p ps=2.72u w=1u l=0.13u
X53 VDD a_53022_43738# a_53085_40283# VDD sg13_lv_pmos ad=0.104p pd=1.34u as=59.75f ps=0.745u w=0.2u l=0.13u
X54 a_53968_20434# a_53738_20514# a_54324_20259# VSS sg13_lv_nmos ad=79.8f pd=0.8u as=54.6f ps=0.68u w=0.42u l=0.13u
X55 VSS 3bit_freq_divider_0.sg13g2_or3_1_0.B a_51648_21103# VSS sg13_lv_nmos ad=0.1045p pd=0.93u as=0.198p ps=1.27u w=0.55u l=0.13u
X56 VDD 3bit_freq_divider_0.EN charge_pump_0.bias_p VDD sg13_lv_pmos ad=0.17p pd=1.68u as=0.17p ps=1.68u w=0.5u l=0.15u
X57 a_55345_23141# 3bit_freq_divider_0.freq_div_cell_0.Cin a_55485_23233# VSS sg13_lv_nmos ad=0.2176p pd=1.96u as=0.1216p ps=1.02u w=0.64u l=0.13u
X58 charge_pump_0.bias_n charge_pump_0.bias_p a_55862_56737# VDD sg13_lv_pmos ad=0.68p pd=4.68u as=0.38p ps=2.38u w=2u l=1u
X59 a_53152_43159# a_52944_43077# a_53058_43159# VDD sg13_lv_pmos ad=0.1106p pd=0.945u as=0.17p ps=1.68u w=0.5u l=0.13u
X60 VDD a_53022_43738# a_55769_40283# VDD sg13_lv_pmos ad=59f pd=0.74u as=59f ps=0.74u w=0.2u l=0.13u
X61 3bit_freq_divider_1.sg13g2_tiehi_1.L_HI a_60584_24580# a_60385_24558# VDD sg13_lv_pmos ad=0.3927p pd=2.99u as=0.4657p ps=2.54u w=1.155u l=0.13u
X62 a_54324_20259# a_53899_20488# a_54252_20259# VSS sg13_lv_nmos ad=54.6f pd=0.68u as=48.3f ps=0.65u w=0.42u l=0.13u
X63 a_62270_24055# a_62119_24117# VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0.34p ps=2.68u w=1u l=0.13u
X64 a_62324_22016# a_62270_22299# a_62246_22016# VSS sg13_lv_nmos ad=48.3f pd=0.65u as=54.6f ps=0.68u w=0.42u l=0.13u
X65 VDD X2 a_52924_21129# VDD sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X66 a_52944_43077# a_53147_40413# a_53085_40283# VDD sg13_lv_pmos ad=0.11p pd=0.94u as=0.17p ps=1.68u w=0.5u l=0.13u
X67 VSS a_53774_21934# a_53738_22270# VSS sg13_lv_nmos ad=0.1544p pd=1.235u as=0.2516p ps=2.16u w=0.74u l=0.13u
X68 a_46749_30782# CLK_IN a_45579_29803# VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=79.8f ps=0.8u w=0.42u l=0.15u
X69 a_54400_43159# a_53152_43159# a_54494_43159# VDD sg13_lv_pmos ad=0.11p pd=0.94u as=0.1106p ps=0.945u w=0.5u l=0.13u
X70 3bit_freq_divider_1.freq_div_cell_0.Cin a_60967_24990# VDD VDD sg13_lv_pmos ad=0.3808p pd=2.92u as=0.1918p ps=1.5u w=1.12u l=0.13u
X71 a_55742_43159# a_53022_43738# VDD VDD sg13_lv_pmos ad=59.75f pd=0.745u as=0.104p ps=1.34u w=0.2u l=0.13u
X72 a_53968_23946# a_53738_24026# a_54324_23771# VSS sg13_lv_nmos ad=79.8f pd=0.8u as=54.6f ps=0.68u w=0.42u l=0.13u
X73 a_63038_20215# 3bit_freq_divider_1.dff_nclk_0.nCLK VSS VSS sg13_lv_nmos ad=47.25f pd=0.645u as=90.3f ps=0.85u w=0.42u l=0.13u
X74 a_62900_20179# a_62654_20215# a_63038_20215# VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=47.25f ps=0.645u w=0.42u l=0.13u
X75 3bit_freq_divider_0.sg13g2_or3_1_0.C a_52886_24904# VSS VSS sg13_lv_nmos ad=0.1628p pd=1.18u as=0.3108p ps=2.32u w=0.74u l=0.13u
X76 VDD a_53022_43738# a_57111_40283# VDD sg13_lv_pmos ad=59f pd=0.74u as=59f ps=0.74u w=0.2u l=0.13u
X77 a_48909_28913# PFD_0.VCO_CLK a_47954_28913# VSS sg13_lv_nmos ad=0.1224p pd=1.4u as=68.39999f ps=0.74u w=0.36u l=0.15u
X78 a_54324_23771# a_53899_24000# a_54252_23771# VSS sg13_lv_nmos ad=54.6f pd=0.68u as=48.3f ps=0.65u w=0.42u l=0.13u
X79 VSS vco_wob_0.vctl a_58454_40850# VSS sg13_lv_nmos ad=0.102p pd=1.28u as=65.99999f ps=0.74u w=0.3u l=0.13u
X80 a_58453_40283# a_53022_43738# VDD VDD sg13_lv_pmos ad=59f pd=0.74u as=0.104p ps=1.34u w=0.2u l=0.13u
X81 a_53899_22244# a_53774_21934# a_53065_21935# VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0.17695p ps=1.56u w=1u l=0.13u
X82 VDD X0 a_52924_24641# VDD sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X83 VDD a_64384_21091# 3bit_freq_divider_1.dff_nclk_0.nCLK VDD sg13_lv_pmos ad=0.3822p pd=1.84u as=0.3808p ps=2.92u w=1.12u l=0.13u
X84 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.D 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.Q a_61972_23244# VSS sg13_lv_nmos ad=0.1628p pd=1.18u as=88.8f ps=0.98u w=0.74u l=0.13u
X85 VDD 3bit_freq_divider_1.sg13g2_tiehi_1.L_HI a_61878_24642# VDD sg13_lv_pmos ad=0.2128p pd=1.5u as=0.3808p ps=2.92u w=1.12u l=0.13u
X86 3bit_freq_divider_1.sg13g2_or3_1_0.B a_63255_23244# a_63426_22886# VDD sg13_lv_pmos ad=0.3808p pd=2.92u as=0.2128p ps=1.5u w=1.12u l=0.13u
X87 VSS vco_wob_0.vctl a_53022_43738# VSS sg13_lv_nmos ad=0.102p pd=1.28u as=65.99999f ps=0.74u w=0.3u l=0.13u
X88 a_51729_23026# a_51631_22774# a_51693_23426# VDD sg13_lv_pmos ad=51.45f pd=0.665u as=79.8f ps=0.8u w=0.42u l=0.13u
X89 a_53147_40413# VSS cap_cmim l=6.99u w=6.99u
X90 a_57084_43159# a_53022_43738# VDD VDD sg13_lv_pmos ad=59.75f pd=0.745u as=0.104p ps=1.34u w=0.2u l=0.13u
X91 a_61887_20534# a_61691_20534# VSS VSS sg13_lv_nmos ad=0.2516p pd=2.16u as=0.1544p ps=1.235u w=0.74u l=0.13u
X92 a_54400_43159# a_53152_43159# a_54494_43159# VDD sg13_lv_pmos ad=0.17p pd=1.68u as=0.11p ps=0.94u w=0.5u l=0.13u
X93 a_62119_22361# a_61691_22290# a_61394_21976# VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0.1428p ps=1.52u w=0.42u l=0.13u
X94 a_52950_23913# a_53065_23691# VDD VDD sg13_lv_pmos ad=0.2856p pd=2.36u as=0.2016p ps=1.5u w=0.84u l=0.13u
X95 a_54504_20259# a_53738_20514# a_53968_20434# VDD sg13_lv_pmos ad=0.1428p pd=1.52u as=79.8f ps=0.8u w=0.42u l=0.13u
X96 a_62119_24117# 3bit_freq_divider_1.dff_nclk_0.nCLK VDD VDD sg13_lv_pmos ad=0.1533p pd=1.57u as=0.11785p ps=1.025u w=0.42u l=0.13u
X97 PFD_0.VCO_CLK PFD_0.VCO_CLK a_46817_27899# VDD sg13_lv_pmos ad=60.8f pd=0.7u as=0.1088p ps=1.32u w=0.32u l=0.15u
X98 VDD 3bit_freq_divider_0.CLK_IN 3bit_freq_divider_1.sg13g2_nand2_1_0.Y VDD sg13_lv_pmos ad=0.3808p pd=2.92u as=0.2128p ps=1.5u w=1.12u l=0.13u
X99 VDD a_62900_21935# a_62879_22369# VDD sg13_lv_pmos ad=79.8f pd=0.8u as=43.05f ps=0.625u w=0.42u l=0.13u
X100 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 3bit_freq_divider_1.sg13g2_nand2_1_0.Y VDD VDD sg13_lv_pmos ad=0.392p pd=2.94u as=0.392p ps=2.94u w=1.12u l=0.13u
X101 a_53350_21129# X2 a_52886_21392# VDD sg13_lv_pmos ad=0.1225p pd=1.245u as=0.34p ps=2.68u w=1u l=0.13u
X102 a_58454_40850# a_58515_40413# a_57173_40413# VSS sg13_lv_nmos ad=0.17p pd=1.68u as=0.11p ps=0.94u w=0.5u l=0.13u
X103 VSS 3bit_freq_divider_0.EN a_56055_21027# VSS sg13_lv_nmos ad=0.2516p pd=2.16u as=66.6f ps=0.92u w=0.74u l=0.13u
X104 VDD a_62654_23727# a_63463_23728# VDD sg13_lv_pmos ad=0.2016p pd=1.5u as=0.2856p ps=2.36u w=0.84u l=0.13u
X105 VSS charge_pump_0.vout VSS VSS sg13_lv_nmos ad=0.285p pd=1.88u as=0 ps=0 w=1.5u l=0.65u
X106 a_55742_43159# a_54494_43159# a_55836_43159# VDD sg13_lv_pmos ad=0.17p pd=1.68u as=0.11p ps=0.94u w=0.5u l=0.13u
X107 a_62654_21971# a_61887_22290# a_62270_22299# VSS sg13_lv_nmos ad=0.2017p pd=1.48u as=0.19397p ps=1.29u w=0.64u l=0.13u
X108 VSS a_62900_20179# a_62848_20215# VSS sg13_lv_nmos ad=90.3f pd=0.85u as=54.6f ps=0.68u w=0.42u l=0.13u
X109 VSS 3bit_freq_divider_0.sg13g2_nand2_1_0.Y 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK VSS sg13_lv_nmos ad=0.259p pd=2.18u as=0.259p ps=2.18u w=0.74u l=0.13u
X110 a_61394_23732# 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.D VDD VDD sg13_lv_pmos ad=79.8f pd=0.8u as=0.1428p ps=1.52u w=0.42u l=0.13u
X111 a_62848_20215# a_61691_20534# a_62654_20215# VSS sg13_lv_nmos ad=54.6f pd=0.68u as=0.2017p ps=1.48u w=0.42u l=0.13u
X112 a_53774_21934# 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK VSS VSS sg13_lv_nmos ad=0.2516p pd=2.16u as=0.1544p ps=1.235u w=0.74u l=0.13u
X113 a_53054_23243# X1 3bit_freq_divider_0.sg13g2_or3_1_0.B VSS sg13_lv_nmos ad=88.8f pd=0.98u as=0.1628p ps=1.18u w=0.74u l=0.13u
X114 a_53350_24641# X0 a_52886_24904# VDD sg13_lv_pmos ad=0.1225p pd=1.245u as=0.34p ps=2.68u w=1u l=0.13u
X115 VDD a_53022_43738# a_58426_43159# VDD sg13_lv_pmos ad=0.104p pd=1.34u as=59f ps=0.74u w=0.2u l=0.13u
X116 a_56038_24617# a_55941_24882# 3bit_freq_divider_0.sg13g2_tiehi_1.L_HI VDD sg13_lv_pmos ad=0.4657p pd=2.54u as=0.3927p ps=2.99u w=1.155u l=0.13u
X117 VDD 3bit_freq_divider_0.dff_nclk_0.nCLK a_53445_20214# VDD sg13_lv_pmos ad=79.8f pd=0.8u as=79.8f ps=0.8u w=0.42u l=0.13u
X118 VSS charge_pump_0.vout VSS VSS sg13_lv_nmos ad=0.285p pd=1.88u as=0 ps=0 w=1.5u l=0.65u
X119 a_57112_40850# vco_wob_0.vctl VSS VSS sg13_lv_nmos ad=65.99999f pd=0.74u as=0.102p ps=1.28u w=0.3u l=0.13u
X120 a_60584_24580# a_60385_24717# a_60479_25023# VSS sg13_lv_nmos ad=0.27427p pd=2.28u as=0.2307p ps=1.615u w=0.795u l=0.13u
X121 VSS a_61707_21488# 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.D VSS sg13_lv_nmos ad=0.3108p pd=2.32u as=0.1628p ps=1.18u w=0.74u l=0.13u
X122 a_63255_25000# Y0 a_63223_24642# VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0.1225p ps=1.245u w=1u l=0.13u
X123 VDD a_51648_24041# a_51685_23725# VDD sg13_lv_pmos ad=0.2163p pd=1.55u as=79.8f ps=0.8u w=0.42u l=0.13u
X124 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.Q a_63463_20216# VDD VDD sg13_lv_pmos ad=0.3808p pd=2.92u as=0.2016p ps=1.5u w=1.12u l=0.13u
X125 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.D a_54434_21392# VSS VSS sg13_lv_nmos ad=0.1628p pd=1.18u as=0.3108p ps=2.32u w=0.74u l=0.13u
X126 VSS Y0 a_63255_25000# VSS sg13_lv_nmos ad=0.15245p pd=1.17u as=0.17462p ps=1.185u w=0.55u l=0.13u
X127 VSS a_56887_49467# VSS VSS sg13_lv_nmos ad=95f pd=0.88u as=0 ps=0 w=0.5u l=0.65u
X128 a_48909_28913# PFD_0.VCO_CLK a_47954_28913# VSS sg13_lv_nmos ad=68.39999f pd=0.74u as=0.1224p ps=1.4u w=0.36u l=0.15u
X129 VDD a_62270_20543# a_62221_20605# VDD sg13_lv_pmos ad=0.11785p pd=1.025u as=51.45f ps=0.665u w=0.42u l=0.13u
X130 a_62246_22016# a_61887_22290# a_62119_22361# VSS sg13_lv_nmos ad=54.6f pd=0.68u as=79.8f ps=0.8u w=0.42u l=0.13u
X131 VDD 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.Q a_63426_21130# VDD sg13_lv_pmos ad=0.2128p pd=1.5u as=0.3808p ps=2.92u w=1.12u l=0.13u
X132 VDD 3bit_freq_divider_0.freq_div_cell_0.Cout a_54898_21129# VDD sg13_lv_pmos ad=0.36p pd=2.72u as=0.1225p ps=1.245u w=1u l=0.13u
X133 VSS charge_pump_0.vout VSS VSS sg13_lv_nmos ad=0.285p pd=1.88u as=0 ps=0 w=1.5u l=0.65u
X134 a_64362_24865# a_64459_24995# a_64731_24890# VDD sg13_lv_pmos ad=0.2442p pd=2.06u as=0.4657p ps=2.54u w=0.66u l=0.13u
X135 a_55831_40413# a_57173_40413# a_57112_40850# VSS sg13_lv_nmos ad=0.11p pd=0.94u as=0.17p ps=1.68u w=0.5u l=0.13u
X136 VSS a_56887_49467# VSS VSS sg13_lv_nmos ad=95f pd=0.88u as=0 ps=0 w=0.5u l=0.65u
X137 a_47777_29803# a_46749_30782# VSS VSS sg13_lv_nmos ad=0.1224p pd=1.4u as=0.1224p ps=1.4u w=0.36u l=0.15u
X138 a_55086_21975# 3bit_freq_divider_0.dff_nclk_0.nCLK VSS VSS sg13_lv_nmos ad=50.4f pd=0.66u as=0.1428p ps=1.52u w=0.42u l=0.13u
X139 VDD 3bit_freq_divider_0.sg13g2_tiehi_1.L_HI a_54898_24641# VDD sg13_lv_pmos ad=0.36p pd=2.72u as=0.1225p ps=1.245u w=1u l=0.13u
X140 a_53445_21970# a_53065_21935# VDD VDD sg13_lv_pmos ad=79.8f pd=0.8u as=0.2163p ps=1.55u w=0.42u l=0.13u
X141 VSS 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.Q a_52886_23148# VSS sg13_lv_nmos ad=0.374p pd=2.46u as=0.17462p ps=1.185u w=0.55u l=0.13u
X142 a_64384_21091# 3bit_freq_divider_1.sg13g2_or3_1_0.A VSS VSS sg13_lv_nmos ad=0.198p pd=1.27u as=0.13395p ps=1.12u w=0.55u l=0.13u
X143 a_63255_23244# 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.Q VSS VSS sg13_lv_nmos ad=0.17462p pd=1.185u as=0.374p ps=2.46u w=0.55u l=0.13u
X144 a_54494_43159# a_53152_43159# a_54400_43159# VDD sg13_lv_pmos ad=0.1106p pd=0.945u as=0.17p ps=1.68u w=0.5u l=0.13u
X145 a_63426_24642# Y0 VDD VDD sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X146 a_62270_20543# a_62119_20605# VSS VSS sg13_lv_nmos ad=0.19397p pd=1.29u as=0.1825p ps=1.325u w=0.64u l=0.13u
X147 VSS a_56887_49467# VSS VSS sg13_lv_nmos ad=95f pd=0.88u as=0 ps=0 w=0.5u l=0.65u
X148 VSS vco_wob_0.vctl a_58653_42591# VSS sg13_lv_nmos ad=0.102p pd=1.28u as=65.99999f ps=0.74u w=0.3u l=0.13u
X149 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.nQ a_62654_21971# VSS VSS sg13_lv_nmos ad=0.2775p pd=2.23u as=0.2516p ps=2.16u w=0.74u l=0.13u
X150 a_58653_42591# a_57178_43159# 3bit_freq_divider_0.CLK_IN VSS sg13_lv_nmos ad=0.17p pd=1.68u as=0.11p ps=0.94u w=0.5u l=0.13u
X151 VDD a_64383_23889# a_64384_24445# VDD sg13_lv_pmos ad=0.2016p pd=1.5u as=0.2856p ps=2.36u w=0.84u l=0.13u
X152 a_51708_21299# 3bit_freq_divider_0.sg13g2_or3_1_0.A VDD VDD sg13_lv_pmos ad=0.22p pd=1.44u as=0.3822p ps=1.84u w=1u l=0.13u
X153 VSS 3bit_freq_divider_0.dff_nclk_0.nRST a_52074_23129# VSS sg13_lv_nmos ad=0.1825p pd=1.325u as=48.3f ps=0.65u w=0.42u l=0.13u
X154 a_53147_40413# a_54489_40413# a_54427_40283# VDD sg13_lv_pmos ad=0.11p pd=0.94u as=0.17p ps=1.68u w=0.5u l=0.13u
X155 VDD 3bit_freq_divider_0.sg13g2_nand2_1_0.Y 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.sg13g2_dfrbp_1_0.CLK VDD sg13_lv_pmos ad=0.392p pd=2.94u as=0.392p ps=2.94u w=1.12u l=0.13u
X156 a_57178_43159# VSS cap_cmim l=6.99u w=6.99u
X157 VSS charge_pump_0.vout VSS VSS sg13_lv_nmos ad=0.51p pd=3.68u as=0 ps=0 w=1.5u l=0.65u
X158 VSS charge_pump_0.vout VSS VSS sg13_lv_nmos ad=0.285p pd=1.88u as=0 ps=0 w=1.5u l=0.65u
X159 VSS a_56887_49467# VSS VSS sg13_lv_nmos ad=95f pd=0.88u as=0 ps=0 w=0.5u l=0.65u
X160 a_62879_20613# a_61887_20534# a_62654_20215# VDD sg13_lv_pmos ad=43.05f pd=0.625u as=0.17695p ps=1.56u w=0.42u l=0.13u
X161 a_61887_22290# a_61691_22290# VSS VSS sg13_lv_nmos ad=0.2516p pd=2.16u as=0.1544p ps=1.235u w=0.74u l=0.13u
X162 VSS a_52950_22157# 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.Q VSS sg13_lv_nmos ad=0.14505p pd=1.15u as=0.2516p ps=2.16u w=0.74u l=0.13u
X163 VSS a_56887_49467# VSS VSS sg13_lv_nmos ad=95f pd=0.88u as=0 ps=0 w=0.5u l=0.65u
X164 a_63520_25000# 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.Q VSS VSS sg13_lv_nmos ad=88.8f pd=0.98u as=0.15245p ps=1.17u w=0.74u l=0.13u
X165 a_53702_24124# a_53445_23726# VDD VDD sg13_lv_pmos ad=43.05f pd=0.625u as=79.8f ps=0.8u w=0.42u l=0.13u
X166 a_61707_25000# 3bit_freq_divider_1.sg13g2_tiehi_1.L_HI VSS VSS sg13_lv_nmos ad=0.17462p pd=1.185u as=0.374p ps=2.46u w=0.55u l=0.13u
X167 VDD 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK a_61691_22290# VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0.34p ps=2.68u w=1u l=0.13u
X168 VDD 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.Q a_54472_21129# VDD sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X169 VSS 3bit_freq_divider_0.freq_div_cell_0.Cin a_54602_23243# VSS sg13_lv_nmos ad=0.15245p pd=1.17u as=88.8f ps=0.98u w=0.74u l=0.13u
X170 VSS a_51648_24041# a_51648_24438# VSS sg13_lv_nmos ad=0.14505p pd=1.15u as=0.187p ps=1.78u w=0.55u l=0.13u
X171 VSS charge_pump_0.vout VSS VSS sg13_lv_nmos ad=0.285p pd=1.88u as=0 ps=0 w=1.5u l=0.65u
X172 a_53147_40413# a_54489_40413# a_54427_40283# VDD sg13_lv_pmos ad=0.1106p pd=0.945u as=0.11p ps=0.94u w=0.5u l=0.13u
X173 a_62270_20543# a_62119_20605# VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0.34p ps=2.68u w=1u l=0.13u
X174 a_51648_21103# 3bit_freq_divider_0.sg13g2_or3_1_0.C a_51708_21413# VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0.1275p ps=1.255u w=1u l=0.13u
X175 VDD 3bit_freq_divider_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK a_51631_22774# VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0.34p ps=2.68u w=1u l=0.13u
X176 VSS vco_wob_0.vctl a_53086_40850# VSS sg13_lv_nmos ad=0.102p pd=1.28u as=65.99999f ps=0.74u w=0.3u l=0.13u
X177 a_59800_40852# vco_wob_0.vctl VSS VSS sg13_lv_nmos ad=65.99999f pd=0.74u as=0.102p ps=1.28u w=0.3u l=0.13u
X178 VSS a_56887_49467# VSS VSS sg13_lv_nmos ad=95f pd=0.88u as=0 ps=0 w=0.5u l=0.65u
X179 a_53085_40283# a_53022_43738# VDD VDD sg13_lv_pmos ad=59f pd=0.74u as=0.104p ps=1.34u w=0.2u l=0.13u
X180 a_62654_23727# a_61887_24046# a_62270_24055# VSS sg13_lv_nmos ad=0.2017p pd=1.48u as=0.19397p ps=1.29u w=0.64u l=0.13u
X181 3bit_freq_divider_0.EN nEN VDD VDD sg13_lv_pmos ad=0.392p pd=2.94u as=0.392p ps=2.94u w=1.12u l=0.13u
X182 VDD a_58734_56203# a_58734_56203# VDD sg13_lv_pmos ad=0.17p pd=1.68u as=0.17p ps=1.68u w=0.5u l=0.15u
X183 VDD a_64383_23706# a_64817_23685# VDD sg13_lv_pmos ad=79.8f pd=0.8u as=43.05f ps=0.625u w=0.42u l=0.13u
X184 VDD 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.Q a_54472_24641# VDD sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X185 VSS 3bit_freq_divider_0.sg13g2_nand2_1_0.Y 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.sg13g2_dfrbp_1_0.CLK VSS sg13_lv_nmos ad=0.259p pd=2.18u as=0.259p ps=2.18u w=0.74u l=0.13u
X186 a_55862_56737# VDD rhigh l=12u w=1u
X187 VDD a_46817_27899# a_45658_27900# VDD sg13_lv_pmos ad=0.1224p pd=1.4u as=68.39999f ps=0.74u w=0.36u l=0.15u
X188 3bit_freq_divider_1.sg13g2_or3_1_0.B Y1 a_63520_23244# VSS sg13_lv_nmos ad=0.1628p pd=1.18u as=88.8f ps=0.98u w=0.74u l=0.13u
X189 VSS charge_pump_0.vout VSS VSS sg13_lv_nmos ad=0.285p pd=1.88u as=0 ps=0 w=1.5u l=0.65u
X190 a_54489_40413# a_55831_40413# a_55769_40283# VDD sg13_lv_pmos ad=0.1106p pd=0.945u as=0.11p ps=0.94u w=0.5u l=0.13u
X191 a_57084_43159# a_55836_43159# a_57178_43159# VDD sg13_lv_pmos ad=0.17p pd=1.68u as=0.11p ps=0.94u w=0.5u l=0.13u
X192 a_63223_24642# 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.Q VDD VDD sg13_lv_pmos ad=0.1225p pd=1.245u as=0.36p ps=2.72u w=1u l=0.13u
X193 3bit_freq_divider_0.CLK_IN a_57178_43159# a_58426_43159# VDD sg13_lv_pmos ad=0.11p pd=0.94u as=0.11p ps=0.94u w=0.5u l=0.13u
X194 a_58515_40413# 3bit_freq_divider_0.CLK_IN a_59800_40852# VSS sg13_lv_nmos ad=0.11p pd=0.94u as=0.17p ps=1.68u w=0.5u l=0.13u
X195 VDD a_62654_20215# a_62900_20179# VDD sg13_lv_pmos ad=0.2163p pd=1.55u as=79.8f ps=0.8u w=0.42u l=0.13u
X196 a_53086_40850# a_53147_40413# a_52944_43077# VSS sg13_lv_nmos ad=0.17p pd=1.68u as=0.11p ps=0.94u w=0.5u l=0.13u
X197 a_64424_22294# 3bit_freq_divider_1.dff_nclk_0.D a_64424_22200# VSS sg13_lv_nmos ad=50.4f pd=0.66u as=0.1428p ps=1.52u w=0.42u l=0.13u
X198 a_61488_23732# 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.D a_61394_23732# VSS sg13_lv_nmos ad=50.4f pd=0.66u as=0.1428p ps=1.52u w=0.42u l=0.13u
X199 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 3bit_freq_divider_1.sg13g2_nand2_1_0.Y VSS VSS sg13_lv_nmos ad=0.259p pd=2.18u as=0.259p ps=2.18u w=0.74u l=0.13u
X200 a_61061_21478# 3bit_freq_divider_1.freq_div_cell_0.Cout a_60967_21478# VSS sg13_lv_nmos ad=0.1216p pd=1.02u as=0.2176p ps=1.96u w=0.64u l=0.13u
X201 VSS 3bit_freq_divider_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK a_51631_22774# VSS sg13_lv_nmos ad=0.1544p pd=1.235u as=0.2516p ps=2.16u w=0.74u l=0.13u
X202 a_62221_20605# a_61691_20534# a_62119_20605# VDD sg13_lv_pmos ad=51.45f pd=0.665u as=79.8f ps=0.8u w=0.42u l=0.13u
X203 VDD a_53022_43738# a_54427_40283# VDD sg13_lv_pmos ad=0.104p pd=1.34u as=59.75f ps=0.745u w=0.2u l=0.13u
X204 VSS a_53968_22190# a_53899_22244# VSS sg13_lv_nmos ad=0.1825p pd=1.325u as=0.19397p ps=1.29u w=0.64u l=0.13u
X205 VSS charge_pump_0.vout VSS VSS sg13_lv_nmos ad=0.285p pd=1.88u as=0 ps=0 w=1.5u l=0.65u
X206 3bit_freq_divider_1.sg13g2_nand2_1_0.Y 3bit_freq_divider_0.CLK_IN a_60531_21028# VSS sg13_lv_nmos ad=0.2516p pd=2.16u as=66.6f ps=0.92u w=0.74u l=0.13u
X207 VSS a_55345_21385# 3bit_freq_divider_0.freq_div_cell_1.Cout VSS sg13_lv_nmos ad=0.1331p pd=1.12u as=0.2516p ps=2.16u w=0.74u l=0.13u
X208 a_59097_54704# 3bit_freq_divider_0.EN VSS VSS sg13_lv_nmos ad=0.17p pd=1.68u as=0.17p ps=1.68u w=0.5u l=0.15u
X209 a_52114_22293# 3bit_freq_divider_0.dff_nclk_0.D a_51684_22284# VSS sg13_lv_nmos ad=50.4f pd=0.66u as=0.1428p ps=1.52u w=0.42u l=0.13u
X210 a_51693_23075# a_51693_23426# VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0.34p ps=2.68u w=1u l=0.13u
X211 VDD a_64383_23889# a_64383_23706# VDD sg13_lv_pmos ad=0.2163p pd=1.55u as=79.8f ps=0.8u w=0.42u l=0.13u
X212 a_61061_24990# 3bit_freq_divider_1.sg13g2_tiehi_1.L_HI a_60967_24990# VSS sg13_lv_nmos ad=0.1216p pd=1.02u as=0.2176p ps=1.96u w=0.64u l=0.13u
X213 a_58515_40413# VSS cap_cmim l=6.99u w=6.99u
X214 a_54472_21129# 3bit_freq_divider_0.freq_div_cell_0.Cout VDD VDD sg13_lv_pmos ad=0.3808p pd=2.92u as=0.2128p ps=1.5u w=1.12u l=0.13u
X215 a_61887_22290# a_61691_22290# VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0.19p ps=1.38u w=1u l=0.13u
X216 VDD a_53022_43738# a_53058_43159# VDD sg13_lv_pmos ad=0.104p pd=1.34u as=59f ps=0.74u w=0.2u l=0.13u
X217 a_61878_24642# 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.Q VDD VDD sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X218 VSS 3bit_freq_divider_1.dff_nclk_0.nCLK a_61488_21976# VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=50.4f ps=0.66u w=0.42u l=0.13u
X219 a_54400_43159# a_53022_43738# VDD VDD sg13_lv_pmos ad=59f pd=0.74u as=59f ps=0.74u w=0.2u l=0.13u
X220 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.Q a_63463_20216# VSS VSS sg13_lv_nmos ad=0.2516p pd=2.16u as=0.14505p ps=1.15u w=0.74u l=0.13u
X221 a_54434_23148# 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.Q VSS VSS sg13_lv_nmos ad=0.17462p pd=1.185u as=0.15245p ps=1.17u w=0.55u l=0.13u
X222 VDD a_53022_43738# a_55769_40283# VDD sg13_lv_pmos ad=0.104p pd=1.34u as=59.75f ps=0.745u w=0.2u l=0.13u
X223 3bit_freq_divider_0.dff_nclk_0.D a_51648_24041# VDD VDD sg13_lv_pmos ad=0.7616p pd=3.6u as=0.2163p ps=1.55u w=1.12u l=0.13u
X224 3bit_freq_divider_1.freq_div_cell_0.Cout a_60967_23234# VSS VSS sg13_lv_nmos ad=0.2516p pd=2.16u as=0.1331p ps=1.12u w=0.74u l=0.13u
X225 VSS a_56887_49467# VSS VSS sg13_lv_nmos ad=95f pd=0.88u as=0 ps=0 w=0.5u l=0.65u
X226 a_54472_24641# 3bit_freq_divider_0.sg13g2_tiehi_1.L_HI VDD VDD sg13_lv_pmos ad=0.3808p pd=2.92u as=0.2128p ps=1.5u w=1.12u l=0.13u
X227 a_55485_24989# 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.Q VSS VSS sg13_lv_nmos ad=0.1216p pd=1.02u as=0.1331p ps=1.12u w=0.64u l=0.13u
X228 PFD_0.VCO_CLK a_51648_24438# VSS VSS sg13_lv_nmos ad=0.2516p pd=2.16u as=0.14505p ps=1.15u w=0.74u l=0.13u
X229 a_62900_21935# 3bit_freq_divider_1.dff_nclk_0.nCLK VDD VDD sg13_lv_pmos ad=79.8f pd=0.8u as=79.8f ps=0.8u w=0.42u l=0.13u
X230 a_53774_21934# 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0.19p ps=1.38u w=1u l=0.13u
X231 a_55742_43159# a_53022_43738# VDD VDD sg13_lv_pmos ad=59f pd=0.74u as=59f ps=0.74u w=0.2u l=0.13u
X232 a_53899_22244# a_53738_22270# a_53065_21935# VSS sg13_lv_nmos ad=0.19397p pd=1.29u as=0.2017p ps=1.48u w=0.64u l=0.13u
X233 a_64383_23889# a_64383_23628# a_64419_23326# VDD sg13_lv_pmos ad=0.17695p pd=1.56u as=0.19p ps=1.38u w=1u l=0.13u
X234 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.nQ a_62654_23727# VSS VSS sg13_lv_nmos ad=0.2775p pd=2.23u as=0.2516p ps=2.16u w=0.74u l=0.13u
X235 3bit_freq_divider_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 3bit_freq_divider_0.dff_nclk_0.nCLK VDD VDD sg13_lv_pmos ad=0.392p pd=2.94u as=0.392p ps=2.94u w=1.12u l=0.13u
X236 a_58426_43159# a_53022_43738# VDD VDD sg13_lv_pmos ad=59.75f pd=0.745u as=0.104p ps=1.34u w=0.2u l=0.13u
X237 VSS 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.Q a_53054_23243# VSS sg13_lv_nmos ad=0.15245p pd=1.17u as=88.8f ps=0.98u w=0.74u l=0.13u
X238 VSS Y2 a_63255_21488# VSS sg13_lv_nmos ad=0.15245p pd=1.17u as=0.17462p ps=1.185u w=0.55u l=0.13u
X239 VSS a_56887_49467# VSS VSS sg13_lv_nmos ad=95f pd=0.88u as=0 ps=0 w=0.5u l=0.65u
X240 a_52950_20401# a_53065_20179# VDD VDD sg13_lv_pmos ad=0.2856p pd=2.36u as=0.2016p ps=1.5u w=0.84u l=0.13u
X241 a_62119_20605# 3bit_freq_divider_1.dff_nclk_0.nCLK VDD VDD sg13_lv_pmos ad=0.1533p pd=1.57u as=0.11785p ps=1.025u w=0.42u l=0.13u
X242 a_60531_21028# 3bit_freq_divider_0.EN VSS VSS sg13_lv_nmos ad=66.6f pd=0.92u as=0.2516p ps=2.16u w=0.74u l=0.13u
X243 VDD a_52950_20401# 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.Q VDD sg13_lv_pmos ad=0.2016p pd=1.5u as=0.3808p ps=2.92u w=1.12u l=0.13u
X244 a_47777_29803# a_46749_30782# VDD VDD sg13_lv_pmos ad=0.1224p pd=1.4u as=68.39999f ps=0.74u w=0.36u l=0.15u
X245 VSS a_52950_23913# 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.Q VSS sg13_lv_nmos ad=0.14505p pd=1.15u as=0.2516p ps=2.16u w=0.74u l=0.13u
X246 a_51693_23075# a_51693_23426# VSS VSS sg13_lv_nmos ad=0.19397p pd=1.29u as=0.1825p ps=1.325u w=0.64u l=0.13u
X247 VDD 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.sg13g2_dfrbp_1_0.CLK a_61691_24046# VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0.34p ps=2.68u w=1u l=0.13u
X248 a_54602_24999# 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.Q 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.D VSS sg13_lv_nmos ad=88.8f pd=0.98u as=0.1628p ps=1.18u w=0.74u l=0.13u
X249 a_53065_21935# a_53738_22270# a_53702_22368# VDD sg13_lv_pmos ad=0.17695p pd=1.56u as=43.05f ps=0.625u w=0.42u l=0.13u
X250 VSS vco_wob_0.vctl a_53285_42591# VSS sg13_lv_nmos ad=0.102p pd=1.28u as=65.99999f ps=0.74u w=0.3u l=0.13u
X251 VDD a_62654_20215# a_63463_20216# VDD sg13_lv_pmos ad=0.2016p pd=1.5u as=0.2856p ps=2.36u w=0.84u l=0.13u
X252 a_53285_42591# a_52944_43077# a_53152_43159# VSS sg13_lv_nmos ad=0.17p pd=1.68u as=0.11p ps=0.94u w=0.5u l=0.13u
X253 VDD 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.Q a_60967_23234# VDD sg13_lv_pmos ad=0.1918p pd=1.5u as=0.1596p ps=1.22u w=0.84u l=0.13u
X254 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.D a_61707_25000# a_61878_24642# VDD sg13_lv_pmos ad=0.3808p pd=2.92u as=0.2128p ps=1.5u w=1.12u l=0.13u
X255 3bit_freq_divider_1.freq_div_cell_1.Cout a_60967_21478# VDD VDD sg13_lv_pmos ad=0.3808p pd=2.92u as=0.1918p ps=1.5u w=1.12u l=0.13u
X256 a_54842_49733# a_54357_49278# charge_pump_0.vout VDD sg13_lv_pmos ad=55.5f pd=0.74u as=0.1005p ps=1.34u w=0.15u l=0.13u
X257 a_54494_43159# VSS cap_cmim l=6.99u w=6.99u
X258 a_61707_25000# 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.Q a_61675_24642# VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0.1225p ps=1.245u w=1u l=0.13u
X259 a_61394_20220# 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.D VDD VDD sg13_lv_pmos ad=79.8f pd=0.8u as=0.1428p ps=1.52u w=0.42u l=0.13u
X260 VDD 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.D a_54504_22015# VDD sg13_lv_pmos ad=0.1428p pd=1.52u as=79.8f ps=0.8u w=0.42u l=0.13u
X261 a_55345_23141# 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.Q VDD VDD sg13_lv_pmos ad=0.1596p pd=1.22u as=0.1918p ps=1.5u w=0.84u l=0.13u
X262 charge_pump_0.bias_n nEN VSS VSS sg13_lv_nmos ad=0.17p pd=1.68u as=0.17p ps=1.68u w=0.5u l=0.15u
X263 a_53022_43738# a_53022_43738# VDD VDD sg13_lv_pmos ad=59.75f pd=0.745u as=59f ps=0.74u w=0.2u l=0.13u
X264 VSS 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.Q a_61707_25000# VSS sg13_lv_nmos ad=0.15245p pd=1.17u as=0.17462p ps=1.185u w=0.55u l=0.13u
X265 3bit_freq_divider_0.sg13g2_or3_1_0.A a_52886_21392# VSS VSS sg13_lv_nmos ad=0.1628p pd=1.18u as=0.3108p ps=2.32u w=0.74u l=0.13u
X266 VSS charge_pump_0.vout VSS VSS sg13_lv_nmos ad=0.285p pd=1.88u as=0 ps=0 w=1.5u l=0.65u
X267 VSS a_56887_49467# VSS VSS sg13_lv_nmos ad=95f pd=0.88u as=0 ps=0 w=0.5u l=0.65u
X268 a_54427_40283# a_54489_40413# a_53147_40413# VDD sg13_lv_pmos ad=0.17p pd=1.68u as=0.1106p ps=0.945u w=0.5u l=0.13u
X269 a_54252_20259# 3bit_freq_divider_0.dff_nclk_0.nCLK VSS VSS sg13_lv_nmos ad=48.3f pd=0.65u as=0.1825p ps=1.325u w=0.42u l=0.13u
X270 a_54427_40283# a_53022_43738# VDD VDD sg13_lv_pmos ad=59f pd=0.74u as=0.104p ps=1.34u w=0.2u l=0.13u
X271 a_55345_24897# 3bit_freq_divider_0.sg13g2_tiehi_1.L_HI a_55485_24989# VSS sg13_lv_nmos ad=0.2176p pd=1.96u as=0.1216p ps=1.02u w=0.64u l=0.13u
X272 CLK_OUT a_64384_24445# VSS VSS sg13_lv_nmos ad=0.2516p pd=2.16u as=0.14505p ps=1.15u w=0.74u l=0.13u
X273 a_54504_20259# a_53774_20178# a_53968_20434# VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=79.8f ps=0.8u w=0.42u l=0.13u
X274 VSS charge_pump_0.vout VSS VSS sg13_lv_nmos ad=0.285p pd=1.88u as=0 ps=0 w=1.5u l=0.65u
X275 VSS a_51685_23725# a_52119_23653# VSS sg13_lv_nmos ad=90.3f pd=0.85u as=54.6f ps=0.68u w=0.42u l=0.13u
X276 VDD 3bit_freq_divider_1.freq_div_cell_0.Cout a_61878_21130# VDD sg13_lv_pmos ad=0.2128p pd=1.5u as=0.3808p ps=2.92u w=1.12u l=0.13u
X277 a_52950_22157# a_53065_21935# VSS VSS sg13_lv_nmos ad=0.187p pd=1.78u as=0.14505p ps=1.15u w=0.55u l=0.13u
X278 a_55969_42591# vco_wob_0.vctl VSS VSS sg13_lv_nmos ad=65.99999f pd=0.74u as=0.102p ps=1.28u w=0.3u l=0.13u
X279 a_55836_43159# a_54494_43159# a_55969_42591# VSS sg13_lv_nmos ad=0.11p pd=0.94u as=0.17p ps=1.68u w=0.5u l=0.13u
X280 a_55770_40850# vco_wob_0.vctl VSS VSS sg13_lv_nmos ad=65.99999f pd=0.74u as=0.102p ps=1.28u w=0.3u l=0.13u
X281 a_62654_23727# a_61691_24046# a_62270_24055# VDD sg13_lv_pmos ad=0.17695p pd=1.56u as=0.19p ps=1.38u w=1u l=0.13u
X282 a_64714_21414# 3bit_freq_divider_1.sg13g2_or3_1_0.B a_64714_21300# VDD sg13_lv_pmos ad=0.1275p pd=1.255u as=0.22p ps=1.44u w=1u l=0.13u
X283 VDD a_51648_24041# a_51648_24438# VDD sg13_lv_pmos ad=0.2016p pd=1.5u as=0.2856p ps=2.36u w=0.84u l=0.13u
X284 VSS a_56887_49467# VSS VSS sg13_lv_nmos ad=95f pd=0.88u as=0 ps=0 w=0.5u l=0.65u
X285 a_55831_40413# VSS cap_cmim l=6.99u w=6.99u
X286 a_52924_21129# 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.Q VDD VDD sg13_lv_pmos ad=0.3808p pd=2.92u as=0.2128p ps=1.5u w=1.12u l=0.13u
X287 VSS a_56887_49467# VSS VSS sg13_lv_nmos ad=95f pd=0.88u as=0 ps=0 w=0.5u l=0.65u
X288 a_55769_40283# a_55831_40413# a_54489_40413# VDD sg13_lv_pmos ad=0.17p pd=1.68u as=0.1106p ps=0.945u w=0.5u l=0.13u
X289 VSS a_62654_21971# a_63463_21972# VSS sg13_lv_nmos ad=0.14505p pd=1.15u as=0.187p ps=1.78u w=0.55u l=0.13u
X290 a_54252_23771# 3bit_freq_divider_0.dff_nclk_0.nCLK VSS VSS sg13_lv_nmos ad=48.3f pd=0.65u as=0.1825p ps=1.325u w=0.42u l=0.13u
X291 VDD a_45658_27900# PFD_0.DOWN VDD sg13_lv_pmos ad=0.1088p pd=1.32u as=60.8f ps=0.7u w=0.32u l=0.15u
X292 3bit_freq_divider_1.dff_nclk_0.D a_64383_23889# VDD VDD sg13_lv_pmos ad=0.7616p pd=3.6u as=0.2163p ps=1.55u w=1.12u l=0.13u
X293 a_45658_27900# a_46817_27899# VDD VDD sg13_lv_pmos ad=68.39999f pd=0.74u as=0.1224p ps=1.4u w=0.36u l=0.15u
X294 VSS 3bit_freq_divider_0.dff_nclk_0.nCLK a_53539_21970# VSS sg13_lv_nmos ad=90.3f pd=0.85u as=47.25f ps=0.645u w=0.42u l=0.13u
X295 a_53539_21970# a_53065_21935# a_53445_21970# VSS sg13_lv_nmos ad=47.25f pd=0.645u as=0.1428p ps=1.52u w=0.42u l=0.13u
X296 VDD 3bit_freq_divider_0.dff_nclk_0.nCLK a_53968_22190# VDD sg13_lv_pmos ad=0.11785p pd=1.025u as=0.1533p ps=1.57u w=0.42u l=0.13u
X297 a_54504_23771# a_53774_23690# a_53968_23946# VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=79.8f ps=0.8u w=0.42u l=0.13u
X298 VSS a_53968_23946# a_53899_24000# VSS sg13_lv_nmos ad=0.1825p pd=1.325u as=0.19397p ps=1.29u w=0.64u l=0.13u
X299 a_52924_22885# a_52886_23148# 3bit_freq_divider_0.sg13g2_or3_1_0.B VDD sg13_lv_pmos ad=0.2128p pd=1.5u as=0.3808p ps=2.92u w=1.12u l=0.13u
X300 a_52886_23148# X1 VSS VSS sg13_lv_nmos ad=0.17462p pd=1.185u as=0.15245p ps=1.17u w=0.55u l=0.13u
X301 a_58453_40283# a_58515_40413# a_57173_40413# VDD sg13_lv_pmos ad=0.11p pd=0.94u as=0.11p ps=0.94u w=0.5u l=0.13u
X302 a_63520_21488# 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.Q VSS VSS sg13_lv_nmos ad=88.8f pd=0.98u as=0.15245p ps=1.17u w=0.74u l=0.13u
X303 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.nQ a_62654_23727# VDD VDD sg13_lv_pmos ad=0.7616p pd=3.6u as=0.2163p ps=1.55u w=1.12u l=0.13u
X304 a_54427_40283# a_53022_43738# VDD VDD sg13_lv_pmos ad=59.75f pd=0.745u as=59f ps=0.74u w=0.2u l=0.13u
X305 a_64731_24890# a_64398_24796# 3bit_freq_divider_1.dff_nclk_0.nRST VDD sg13_lv_pmos ad=0.4657p pd=2.54u as=0.3927p ps=2.99u w=1.155u l=0.13u
X306 a_61707_21488# 3bit_freq_divider_1.freq_div_cell_0.Cout VSS VSS sg13_lv_nmos ad=0.17462p pd=1.185u as=0.374p ps=2.46u w=0.55u l=0.13u
X307 VDD a_53968_22190# a_53899_22244# VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0.19p ps=1.38u w=1u l=0.13u
X308 VSS a_56887_49467# VSS VSS sg13_lv_nmos ad=95f pd=0.88u as=0 ps=0 w=0.5u l=0.65u
X309 a_52924_24641# 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.Q VDD VDD sg13_lv_pmos ad=0.3808p pd=2.92u as=0.2128p ps=1.5u w=1.12u l=0.13u
X310 VSS a_56887_49467# VSS VSS sg13_lv_nmos ad=95f pd=0.88u as=0 ps=0 w=0.5u l=0.65u
X311 a_54489_40413# a_55831_40413# a_55770_40850# VSS sg13_lv_nmos ad=0.11p pd=0.94u as=0.17p ps=1.68u w=0.5u l=0.13u
X312 VDD a_52950_23913# 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.Q VDD sg13_lv_pmos ad=0.2016p pd=1.5u as=0.3808p ps=2.92u w=1.12u l=0.13u
X313 a_61887_24046# a_61691_24046# VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0.19p ps=1.38u w=1u l=0.13u
X314 charge_pump_0.vout vco_wob_0.vctl rhigh l=0.96u w=0.6u
X315 VDD a_53065_21935# 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.nQ VDD sg13_lv_pmos ad=0.2163p pd=1.55u as=0.7616p ps=3.6u w=1.12u l=0.13u
X316 a_53152_43159# a_52944_43077# a_53058_43159# VDD sg13_lv_pmos ad=0.11p pd=0.94u as=0.11p ps=0.94u w=0.5u l=0.13u
X317 VDD a_51685_23725# a_51721_23684# VDD sg13_lv_pmos ad=79.8f pd=0.8u as=43.05f ps=0.625u w=0.42u l=0.13u
X318 VDD a_53774_23690# a_53738_24026# VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0.34p ps=2.68u w=1u l=0.13u
X319 a_55836_43159# a_54494_43159# a_55742_43159# VDD sg13_lv_pmos ad=0.1106p pd=0.945u as=0.17p ps=1.68u w=0.5u l=0.13u
X320 a_55769_40283# a_53022_43738# VDD VDD sg13_lv_pmos ad=59.75f pd=0.745u as=59f ps=0.74u w=0.2u l=0.13u
X321 a_56013_24979# a_56137_24678# a_56038_24617# VDD sg13_lv_pmos ad=0.2442p pd=2.06u as=0.4657p ps=2.54u w=0.66u l=0.13u
X322 VDD 3bit_freq_divider_0.freq_div_cell_0.Cin a_55345_23141# VDD sg13_lv_pmos ad=0.2856p pd=2.36u as=0.1596p ps=1.22u w=0.84u l=0.13u
X323 VSS a_56887_49467# VSS VSS sg13_lv_nmos ad=95f pd=0.88u as=0 ps=0 w=0.5u l=0.65u
X324 a_48909_28913# CLK_IN VSS VSS sg13_lv_nmos ad=0.1224p pd=1.4u as=0.1224p ps=1.4u w=0.36u l=0.15u
X325 a_64464_23052# a_64383_23434# a_64383_23300# VSS sg13_lv_nmos ad=54.6f pd=0.68u as=79.8f ps=0.8u w=0.42u l=0.13u
X326 a_56055_21027# 3bit_freq_divider_0.CLK_IN 3bit_freq_divider_0.sg13g2_nand2_1_0.Y VSS sg13_lv_nmos ad=66.6f pd=0.92u as=0.2516p ps=2.16u w=0.74u l=0.13u
X327 VSS a_56887_49467# VSS VSS sg13_lv_nmos ad=95f pd=0.88u as=0 ps=0 w=0.5u l=0.65u
X328 a_61972_25000# 3bit_freq_divider_1.sg13g2_tiehi_1.L_HI VSS VSS sg13_lv_nmos ad=88.8f pd=0.98u as=0.15245p ps=1.17u w=0.74u l=0.13u
X329 a_63255_21488# Y2 a_63223_21130# VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0.1225p ps=1.245u w=1u l=0.13u
X330 a_51648_21103# 3bit_freq_divider_0.sg13g2_or3_1_0.C VSS VSS sg13_lv_nmos ad=0.187p pd=1.78u as=0.1045p ps=0.93u w=0.55u l=0.13u
X331 a_53899_24000# a_53738_24026# a_53065_23691# VSS sg13_lv_nmos ad=0.19397p pd=1.29u as=0.2017p ps=1.48u w=0.64u l=0.13u
X332 VSS 3bit_freq_divider_0.freq_div_cell_0.Cin a_54434_23148# VSS sg13_lv_nmos ad=0.374p pd=2.46u as=0.17462p ps=1.185u w=0.55u l=0.13u
X333 charge_pump_0.vout PFD_0.DOWN a_54747_49259# VSS sg13_lv_nmos ad=0.408p pd=3.08u as=0.207p ps=1.545u w=1.2u l=0.13u
X334 a_52119_23843# 3bit_freq_divider_0.dff_nclk_0.nRST VSS VSS sg13_lv_nmos ad=47.25f pd=0.645u as=90.3f ps=0.85u w=0.42u l=0.13u
X335 PFD_0.UP a_47777_29803# VDD VDD sg13_lv_pmos ad=0.1088p pd=1.32u as=60.8f ps=0.7u w=0.32u l=0.15u
X336 a_53054_24999# X0 3bit_freq_divider_0.sg13g2_or3_1_0.C VSS sg13_lv_nmos ad=88.8f pd=0.98u as=0.1628p ps=1.18u w=0.74u l=0.13u
X337 VSS charge_pump_0.vout VSS VSS sg13_lv_nmos ad=0.285p pd=1.88u as=0 ps=0 w=1.5u l=0.65u
X338 a_57178_43159# a_55836_43159# a_57084_43159# VDD sg13_lv_pmos ad=0.1106p pd=0.945u as=0.17p ps=1.68u w=0.5u l=0.13u
X339 VDD a_55345_21385# 3bit_freq_divider_0.freq_div_cell_1.Cout VDD sg13_lv_pmos ad=0.1918p pd=1.5u as=0.3808p ps=2.92u w=1.12u l=0.13u
X340 VDD 3bit_freq_divider_1.dff_nclk_0.nCLK a_61394_23732# VDD sg13_lv_pmos ad=0.1428p pd=1.52u as=79.8f ps=0.8u w=0.42u l=0.13u
X341 VSS a_56887_49467# VSS VSS sg13_lv_nmos ad=95f pd=0.88u as=0 ps=0 w=0.5u l=0.65u
X342 a_57084_43159# a_53022_43738# VDD VDD sg13_lv_pmos ad=59f pd=0.74u as=59f ps=0.74u w=0.2u l=0.13u
X343 a_53065_21935# a_53774_21934# a_53722_21970# VSS sg13_lv_nmos ad=0.2017p pd=1.48u as=54.6f ps=0.68u w=0.42u l=0.13u
X344 a_53968_22190# a_53774_21934# a_54352_22360# VDD sg13_lv_pmos ad=79.8f pd=0.8u as=51.45f ps=0.665u w=0.42u l=0.13u
X345 a_53702_20612# a_53445_20214# VDD VDD sg13_lv_pmos ad=43.05f pd=0.625u as=79.8f ps=0.8u w=0.42u l=0.13u
X346 VDD a_53022_43738# a_58426_43159# VDD sg13_lv_pmos ad=59f pd=0.74u as=59.75f ps=0.745u w=0.2u l=0.13u
X347 VSS vco_wob_0.vctl a_59800_40852# VSS sg13_lv_nmos ad=0.102p pd=1.28u as=65.99999f ps=0.74u w=0.3u l=0.13u
X348 a_59799_40285# a_53022_43738# VDD VDD sg13_lv_pmos ad=59f pd=0.74u as=0.104p ps=1.34u w=0.2u l=0.13u
X349 a_60967_24990# 3bit_freq_divider_1.sg13g2_tiehi_1.L_HI VDD VDD sg13_lv_pmos ad=0.1596p pd=1.22u as=0.2856p ps=2.36u w=0.84u l=0.13u
X350 VDD a_53022_43738# a_53085_40283# VDD sg13_lv_pmos ad=59f pd=0.74u as=59f ps=0.74u w=0.2u l=0.13u
X351 a_53722_21970# a_53445_21970# VSS VSS sg13_lv_nmos ad=54.6f pd=0.68u as=90.3f ps=0.85u w=0.42u l=0.13u
X352 VSS charge_pump_0.vout VSS VSS sg13_lv_nmos ad=0.285p pd=1.88u as=0 ps=0 w=1.5u l=0.65u
X353 VSS vco_wob_0.vctl a_54428_40850# VSS sg13_lv_nmos ad=0.102p pd=1.28u as=65.99999f ps=0.74u w=0.3u l=0.13u
X354 VSS charge_pump_0.vout VSS VSS sg13_lv_nmos ad=0.285p pd=1.88u as=0 ps=0 w=1.5u l=0.65u
X355 VSS 3bit_freq_divider_1.dff_nclk_0.nCLK a_62324_23772# VSS sg13_lv_nmos ad=0.1825p pd=1.325u as=48.3f ps=0.65u w=0.42u l=0.13u
X356 VDD a_55345_24897# 3bit_freq_divider_0.freq_div_cell_0.Cin VDD sg13_lv_pmos ad=0.1918p pd=1.5u as=0.3808p ps=2.92u w=1.12u l=0.13u
X357 VSS a_63255_23244# 3bit_freq_divider_1.sg13g2_or3_1_0.B VSS sg13_lv_nmos ad=0.3108p pd=2.32u as=0.1628p ps=1.18u w=0.74u l=0.13u
X358 a_61675_24642# 3bit_freq_divider_1.sg13g2_tiehi_1.L_HI VDD VDD sg13_lv_pmos ad=0.1225p pd=1.245u as=0.36p ps=2.72u w=1u l=0.13u
X359 a_53058_43159# a_53022_43738# VDD VDD sg13_lv_pmos ad=59.75f pd=0.745u as=0.104p ps=1.34u w=0.2u l=0.13u
X360 VDD 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.Q a_63426_22886# VDD sg13_lv_pmos ad=0.2128p pd=1.5u as=0.3808p ps=2.92u w=1.12u l=0.13u
X361 3bit_freq_divider_0.sg13g2_nand2_1_0.Y 3bit_freq_divider_0.CLK_IN VDD VDD sg13_lv_pmos ad=0.2128p pd=1.5u as=0.3808p ps=2.92u w=1.12u l=0.13u
X362 a_53968_22190# a_53738_22270# a_54324_22015# VSS sg13_lv_nmos ad=79.8f pd=0.8u as=54.6f ps=0.68u w=0.42u l=0.13u
X363 a_63426_21130# Y2 VDD VDD sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X364 a_57173_40413# VSS cap_cmim l=6.99u w=6.99u
X365 a_61394_21976# 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.D VDD VDD sg13_lv_pmos ad=79.8f pd=0.8u as=0.1428p ps=1.52u w=0.42u l=0.13u
X366 VSS charge_pump_0.vout VSS VSS sg13_lv_nmos ad=0.285p pd=1.88u as=0 ps=0 w=1.5u l=0.65u
X367 a_54324_22015# a_53899_22244# a_54252_22015# VSS sg13_lv_nmos ad=54.6f pd=0.68u as=48.3f ps=0.65u w=0.42u l=0.13u
X368 a_59800_40852# 3bit_freq_divider_0.CLK_IN a_58515_40413# VSS sg13_lv_nmos ad=0.17p pd=1.68u as=0.11p ps=0.94u w=0.5u l=0.13u
X369 a_58734_56203# a_58536_54976# a_58536_54976# VDD sg13_lv_pmos ad=0.17p pd=1.68u as=0.17p ps=1.68u w=0.5u l=0.15u
X370 a_54428_40850# a_54489_40413# a_53147_40413# VSS sg13_lv_nmos ad=0.17p pd=1.68u as=0.11p ps=0.94u w=0.5u l=0.13u
X371 a_52950_23913# a_53065_23691# VSS VSS sg13_lv_nmos ad=0.187p pd=1.78u as=0.14505p ps=1.15u w=0.55u l=0.13u
X372 a_64383_23300# a_64383_23434# a_64424_22200# VDD sg13_lv_pmos ad=79.8f pd=0.8u as=0.1428p ps=1.52u w=0.42u l=0.13u
X373 VSS 3bit_freq_divider_1.sg13g2_or3_1_0.B a_64384_21091# VSS sg13_lv_nmos ad=0.1045p pd=0.93u as=0.198p ps=1.27u w=0.55u l=0.13u
X374 VSS 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.Q a_52886_24904# VSS sg13_lv_nmos ad=0.374p pd=2.46u as=0.17462p ps=1.185u w=0.55u l=0.13u
X375 VDD 3bit_freq_divider_0.dff_nclk_0.nRST a_51684_22284# VDD sg13_lv_pmos ad=0.1428p pd=1.52u as=79.8f ps=0.8u w=0.42u l=0.13u
X376 VDD charge_pump_0.bias_p charge_pump_0.bias_p VDD sg13_lv_pmos ad=0.68p pd=4.68u as=0.68p ps=4.68u w=2u l=1u
X377 a_64459_24995# a_64459_24995# a_64338_24910# VSS sg13_lv_nmos ad=0.102p pd=1.28u as=0.2307p ps=1.615u w=0.3u l=0.13u
X378 VDD 3bit_freq_divider_0.dff_nclk_0.nCLK a_53445_21970# VDD sg13_lv_pmos ad=79.8f pd=0.8u as=79.8f ps=0.8u w=0.42u l=0.13u
X379 VDD PFD_0.UP a_54357_49278# VDD sg13_lv_pmos ad=0.102p pd=1.28u as=0.102p ps=1.28u w=0.3u l=0.13u
X380 VSS a_62654_23727# a_63463_23728# VSS sg13_lv_nmos ad=0.14505p pd=1.15u as=0.187p ps=1.78u w=0.55u l=0.13u
X381 VSS charge_pump_0.vout VSS VSS sg13_lv_nmos ad=0.285p pd=1.88u as=0 ps=0 w=1.5u l=0.65u
X382 a_53899_24000# a_53774_23690# a_53065_23691# VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0.17695p ps=1.56u w=1u l=0.13u
X383 VDD 3bit_freq_divider_0.dff_nclk_0.nCLK a_53968_23946# VDD sg13_lv_pmos ad=0.11785p pd=1.025u as=0.1533p ps=1.57u w=0.42u l=0.13u
X384 a_53539_23726# a_53065_23691# a_53445_23726# VSS sg13_lv_nmos ad=47.25f pd=0.645u as=0.1428p ps=1.52u w=0.42u l=0.13u
X385 VSS 3bit_freq_divider_0.dff_nclk_0.nCLK a_53539_23726# VSS sg13_lv_nmos ad=90.3f pd=0.85u as=47.25f ps=0.645u w=0.42u l=0.13u
X386 a_57311_42591# vco_wob_0.vctl VSS VSS sg13_lv_nmos ad=65.99999f pd=0.74u as=0.102p ps=1.28u w=0.3u l=0.13u
X387 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.D 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.Q a_61972_25000# VSS sg13_lv_nmos ad=0.1628p pd=1.18u as=88.8f ps=0.98u w=0.74u l=0.13u
X388 3bit_freq_divider_1.sg13g2_or3_1_0.C a_63255_25000# a_63426_24642# VDD sg13_lv_pmos ad=0.3808p pd=2.92u as=0.2128p ps=1.5u w=1.12u l=0.13u
X389 a_57178_43159# a_55836_43159# a_57311_42591# VSS sg13_lv_nmos ad=0.11p pd=0.94u as=0.17p ps=1.68u w=0.5u l=0.13u
X390 a_45579_29803# CLK_IN a_45451_28860# VSS sg13_lv_nmos ad=0.1224p pd=1.4u as=68.39999f ps=0.74u w=0.36u l=0.15u
X391 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.Q a_63463_21972# VDD VDD sg13_lv_pmos ad=0.3808p pd=2.92u as=0.2016p ps=1.5u w=1.12u l=0.13u
X392 VSS 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.sg13g2_dfrbp_1_0.CLK a_61691_24046# VSS sg13_lv_nmos ad=0.1544p pd=1.235u as=0.2516p ps=2.16u w=0.74u l=0.13u
X393 VDD 3bit_freq_divider_1.dff_nclk_0.nRST a_64424_22200# VDD sg13_lv_pmos ad=0.1428p pd=1.52u as=79.8f ps=0.8u w=0.42u l=0.13u
X394 VDD a_64419_23326# a_64809_23027# VDD sg13_lv_pmos ad=0.11785p pd=1.025u as=51.45f ps=0.665u w=0.42u l=0.13u
X395 a_64338_24910# a_64362_24865# a_64398_24796# VSS sg13_lv_nmos ad=0.2307p pd=1.615u as=0.27427p ps=2.28u w=0.795u l=0.13u
X396 a_62654_20215# a_61887_20534# a_62270_20543# VSS sg13_lv_nmos ad=0.2017p pd=1.48u as=0.19397p ps=1.29u w=0.64u l=0.13u
X397 PFD_0.DOWN a_45658_27900# VDD VDD sg13_lv_pmos ad=60.8f pd=0.7u as=60.8f ps=0.7u w=0.32u l=0.15u
X398 a_54472_22885# a_54434_23148# 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.D VDD sg13_lv_pmos ad=0.2128p pd=1.5u as=0.3808p ps=2.92u w=1.12u l=0.13u
X399 VDD 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.Q a_53350_22885# VDD sg13_lv_pmos ad=0.36p pd=2.72u as=0.1225p ps=1.245u w=1u l=0.13u
X400 VSS 3bit_freq_divider_0.sg13g2_nand2_1_0.Y 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.sg13g2_dfrbp_1_0.CLK VSS sg13_lv_nmos ad=0.259p pd=2.18u as=0.259p ps=2.18u w=0.74u l=0.13u
X401 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 3bit_freq_divider_1.sg13g2_nand2_1_0.Y VDD VDD sg13_lv_pmos ad=0.392p pd=2.94u as=0.392p ps=2.94u w=1.12u l=0.13u
X402 a_51648_24041# a_51684_22692# a_51693_23075# VSS sg13_lv_nmos ad=0.2017p pd=1.48u as=0.19397p ps=1.29u w=0.64u l=0.13u
X403 VDD a_62900_23691# a_62879_24125# VDD sg13_lv_pmos ad=79.8f pd=0.8u as=43.05f ps=0.625u w=0.42u l=0.13u
X404 VSS 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.Q a_61707_21488# VSS sg13_lv_nmos ad=0.15245p pd=1.17u as=0.17462p ps=1.185u w=0.55u l=0.13u
X405 a_45579_29803# CLK_IN a_45451_28860# VSS sg13_lv_nmos ad=68.39999f pd=0.74u as=68.39999f ps=0.74u w=0.36u l=0.15u
X406 VSS 3bit_freq_divider_1.dff_nclk_0.nRST a_64424_22294# VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=50.4f ps=0.66u w=0.42u l=0.13u
X407 a_45579_29803# CLK_IN VDD VDD sg13_lv_pmos ad=0.1088p pd=1.32u as=60.8f ps=0.7u w=0.32u l=0.15u
X408 VSS 3bit_freq_divider_0.sg13g2_tiehi_1.L_HI a_54602_24999# VSS sg13_lv_nmos ad=0.15245p pd=1.17u as=88.8f ps=0.98u w=0.74u l=0.13u
X409 a_63223_21130# 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.Q VDD VDD sg13_lv_pmos ad=0.1225p pd=1.245u as=0.36p ps=2.72u w=1u l=0.13u
X410 a_58515_40413# 3bit_freq_divider_0.CLK_IN a_59799_40285# VDD sg13_lv_pmos ad=0.11p pd=0.94u as=0.17p ps=1.68u w=0.5u l=0.13u
X411 a_53085_40283# a_53147_40413# a_52944_43077# VDD sg13_lv_pmos ad=0.11p pd=0.94u as=0.11p ps=0.94u w=0.5u l=0.13u
X412 a_58515_40413# 3bit_freq_divider_0.CLK_IN a_59799_40285# VDD sg13_lv_pmos ad=0.1106p pd=0.945u as=0.11p ps=0.94u w=0.5u l=0.13u
X413 a_61488_20220# 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.D a_61394_20220# VSS sg13_lv_nmos ad=50.4f pd=0.66u as=0.1428p ps=1.52u w=0.42u l=0.13u
X414 a_62654_20215# a_61691_20534# a_62270_20543# VDD sg13_lv_pmos ad=0.17695p pd=1.56u as=0.19p ps=1.38u w=1u l=0.13u
X415 a_54494_43159# a_53152_43159# a_54400_43159# VDD sg13_lv_pmos ad=0.11p pd=0.94u as=0.11p ps=0.94u w=0.5u l=0.13u
X416 VSS charge_pump_0.vout VSS VSS sg13_lv_nmos ad=0.285p pd=1.88u as=0 ps=0 w=1.5u l=0.65u
X417 a_55742_43159# a_54494_43159# a_55836_43159# VDD sg13_lv_pmos ad=0.11p pd=0.94u as=0.1106p ps=0.945u w=0.5u l=0.13u
X418 a_46817_27899# PFD_0.VCO_CLK a_47954_28913# VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=79.8f ps=0.8u w=0.42u l=0.15u
X419 VSS 3bit_freq_divider_0.dff_nclk_0.nRST a_52114_22293# VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=50.4f ps=0.66u w=0.42u l=0.13u
X420 VSS a_53065_21935# 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.nQ VSS sg13_lv_nmos ad=0.2516p pd=2.16u as=0.2775p ps=2.23u w=0.74u l=0.13u
X421 VDD a_53022_43738# a_58453_40283# VDD sg13_lv_pmos ad=59f pd=0.74u as=59f ps=0.74u w=0.2u l=0.13u
X422 a_54352_22360# a_53899_22244# VDD VDD sg13_lv_pmos ad=51.45f pd=0.665u as=0.11785p ps=1.025u w=0.42u l=0.13u
X423 VSS a_61707_23244# 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.D VSS sg13_lv_nmos ad=0.3108p pd=2.32u as=0.1628p ps=1.18u w=0.74u l=0.13u
X424 a_54357_49278# PFD_0.UP VSS VSS sg13_lv_nmos ad=0.1005p pd=1.34u as=0.1005p ps=1.34u w=0.15u l=0.13u
X425 a_53968_23946# a_53774_23690# a_54352_24116# VDD sg13_lv_pmos ad=79.8f pd=0.8u as=51.45f ps=0.665u w=0.42u l=0.13u
X426 VDD 3bit_freq_divider_0.sg13g2_nand2_1_0.Y 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK VDD sg13_lv_pmos ad=0.392p pd=2.94u as=0.392p ps=2.94u w=1.12u l=0.13u
X427 VSS a_56887_49467# VSS VSS sg13_lv_nmos ad=0.17p pd=1.68u as=0 ps=0 w=0.5u l=0.65u
X428 a_53065_23691# a_53774_23690# a_53722_23726# VSS sg13_lv_nmos ad=0.2017p pd=1.48u as=54.6f ps=0.68u w=0.42u l=0.13u
X429 a_61878_21130# 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.Q VDD VDD sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X430 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.D a_54434_23148# VSS VSS sg13_lv_nmos ad=0.1628p pd=1.18u as=0.3108p ps=2.32u w=0.74u l=0.13u
X431 VDD 3bit_freq_divider_0.EN a_58536_54976# VDD sg13_lv_pmos ad=0.17p pd=1.68u as=0.17p ps=1.68u w=0.5u l=0.15u
X432 a_57084_43159# a_55836_43159# a_57178_43159# VDD sg13_lv_pmos ad=0.11p pd=0.94u as=0.1106p ps=0.945u w=0.5u l=0.13u
X433 VDD 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.sg13g2_dfrbp_1_0.CLK a_61691_20534# VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0.34p ps=2.68u w=1u l=0.13u
X434 a_53722_23726# a_53445_23726# VSS VSS sg13_lv_nmos ad=54.6f pd=0.68u as=90.3f ps=0.85u w=0.42u l=0.13u
X435 a_55086_20219# 3bit_freq_divider_0.dff_nclk_0.nCLK VSS VSS sg13_lv_nmos ad=50.4f pd=0.66u as=0.1428p ps=1.52u w=0.42u l=0.13u
X436 3bit_freq_divider_0.CLK_IN VSS cap_cmim l=6.99u w=6.99u
X437 3bit_freq_divider_0.CLK_IN a_57178_43159# a_58426_43159# VDD sg13_lv_pmos ad=0.1106p pd=0.945u as=0.17p ps=1.68u w=0.5u l=0.13u
X438 PFD_0.UP a_47777_29803# VDD VDD sg13_lv_pmos ad=60.8f pd=0.7u as=0.1088p ps=1.32u w=0.32u l=0.15u
X439 a_62879_22369# a_61887_22290# a_62654_21971# VDD sg13_lv_pmos ad=43.05f pd=0.625u as=0.17695p ps=1.56u w=0.42u l=0.13u
X440 VDD a_47777_29803# PFD_0.UP VDD sg13_lv_pmos ad=60.8f pd=0.7u as=60.8f ps=0.7u w=0.32u l=0.15u
X441 VSS 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.Q a_61061_21478# VSS sg13_lv_nmos ad=0.1331p pd=1.12u as=0.1216p ps=1.02u w=0.64u l=0.13u
X442 a_51600_24907# a_51622_24863# 3bit_freq_divider_0.dff_nclk_0.nRST VDD sg13_lv_pmos ad=0.4657p pd=2.54u as=0.3927p ps=2.99u w=1.155u l=0.13u
X443 VSS 3bit_freq_divider_1.dff_nclk_0.nRST a_64464_23130# VSS sg13_lv_nmos ad=0.1825p pd=1.325u as=48.3f ps=0.65u w=0.42u l=0.13u
X444 VSS a_56887_49467# VSS VSS sg13_lv_nmos ad=0.17p pd=1.68u as=0 ps=0 w=0.5u l=0.65u
X445 VDD a_46749_30782# a_47777_29803# VDD sg13_lv_pmos ad=68.39999f pd=0.74u as=0.1224p ps=1.4u w=0.36u l=0.15u
X446 a_55485_21477# 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.Q VSS VSS sg13_lv_nmos ad=0.1216p pd=1.02u as=0.1331p ps=1.12u w=0.64u l=0.13u
X447 VSS a_56887_49467# VSS VSS sg13_lv_nmos ad=95f pd=0.88u as=0 ps=0 w=0.5u l=0.65u
X448 VSS vco_wob_0.vctl a_55969_42591# VSS sg13_lv_nmos ad=0.102p pd=1.28u as=65.99999f ps=0.74u w=0.3u l=0.13u
X449 a_55969_42591# a_54494_43159# a_55836_43159# VSS sg13_lv_nmos ad=0.17p pd=1.68u as=0.11p ps=0.94u w=0.5u l=0.13u
X450 VSS vco_wob_0.vctl a_55770_40850# VSS sg13_lv_nmos ad=0.102p pd=1.28u as=65.99999f ps=0.74u w=0.3u l=0.13u
X451 a_53022_43738# vco_wob_0.vctl VSS VSS sg13_lv_nmos ad=65.99999f pd=0.74u as=0.102p ps=1.28u w=0.3u l=0.13u
X452 a_55769_40283# a_53022_43738# VDD VDD sg13_lv_pmos ad=59f pd=0.74u as=0.104p ps=1.34u w=0.2u l=0.13u
X453 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.nQ a_62654_20215# VSS VSS sg13_lv_nmos ad=0.2775p pd=2.23u as=0.2516p ps=2.16u w=0.74u l=0.13u
X454 a_55086_23731# 3bit_freq_divider_0.dff_nclk_0.nCLK VSS VSS sg13_lv_nmos ad=50.4f pd=0.66u as=0.1428p ps=1.52u w=0.42u l=0.13u
X455 VSS 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.Q a_61061_24990# VSS sg13_lv_nmos ad=0.1331p pd=1.12u as=0.1216p ps=1.02u w=0.64u l=0.13u
X456 VSS a_64383_23706# a_64419_23654# VSS sg13_lv_nmos ad=90.3f pd=0.85u as=54.6f ps=0.68u w=0.42u l=0.13u
X457 a_61972_21488# 3bit_freq_divider_1.freq_div_cell_0.Cout VSS VSS sg13_lv_nmos ad=88.8f pd=0.98u as=0.15245p ps=1.17u w=0.74u l=0.13u
X458 VDD a_53022_43738# a_53058_43159# VDD sg13_lv_pmos ad=59f pd=0.74u as=59.75f ps=0.745u w=0.2u l=0.13u
X459 VSS vco_wob_0.vctl VSS VSS sg13_lv_nmos ad=0.1005p pd=1.34u as=0 ps=0 w=0.15u l=0.13u
X460 a_54434_24904# 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.Q VSS VSS sg13_lv_nmos ad=0.17462p pd=1.185u as=0.15245p ps=1.17u w=0.55u l=0.13u
X461 a_53445_23726# a_53065_23691# VDD VDD sg13_lv_pmos ad=79.8f pd=0.8u as=0.2163p ps=1.55u w=0.42u l=0.13u
X462 a_54400_43159# a_53022_43738# VDD VDD sg13_lv_pmos ad=59.75f pd=0.745u as=0.104p ps=1.34u w=0.2u l=0.13u
X463 a_51684_22692# a_51631_22774# VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0.19p ps=1.38u w=1u l=0.13u
X464 VSS a_56887_49467# VSS VSS sg13_lv_nmos ad=95f pd=0.88u as=0 ps=0 w=0.5u l=0.65u
X465 a_57111_40283# a_57173_40413# a_55831_40413# VDD sg13_lv_pmos ad=0.17p pd=1.68u as=0.1106p ps=0.945u w=0.5u l=0.13u
X466 a_63255_25000# 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.Q VSS VSS sg13_lv_nmos ad=0.17462p pd=1.185u as=0.374p ps=2.46u w=0.55u l=0.13u
X467 charge_pump_0.bias_p a_58536_54976# a_59097_54704# VSS sg13_lv_nmos ad=0.17p pd=1.68u as=0.17p ps=1.68u w=0.5u l=0.15u
X468 VSS a_56887_49467# VSS VSS sg13_lv_nmos ad=95f pd=0.88u as=0 ps=0 w=0.5u l=0.65u
X469 3bit_freq_divider_1.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 3bit_freq_divider_1.dff_nclk_0.nCLK VDD VDD sg13_lv_pmos ad=0.392p pd=2.94u as=0.392p ps=2.94u w=1.12u l=0.13u
X470 VSS a_52950_20401# 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.Q VSS sg13_lv_nmos ad=0.14505p pd=1.15u as=0.2516p ps=2.16u w=0.74u l=0.13u
X471 VSS vco_wob_0.vctl a_57112_40850# VSS sg13_lv_nmos ad=0.102p pd=1.28u as=65.99999f ps=0.74u w=0.3u l=0.13u
X472 a_62119_22361# a_61887_22290# a_61394_21976# VDD sg13_lv_pmos ad=79.8f pd=0.8u as=0.1428p ps=1.52u w=0.42u l=0.13u
X473 a_64383_23706# 3bit_freq_divider_1.dff_nclk_0.nRST VDD VDD sg13_lv_pmos ad=79.8f pd=0.8u as=79.8f ps=0.8u w=0.42u l=0.13u
X474 a_57111_40283# a_53022_43738# VDD VDD sg13_lv_pmos ad=59f pd=0.74u as=0.104p ps=1.34u w=0.2u l=0.13u
X475 a_51693_23426# a_51684_22692# a_51684_22284# VDD sg13_lv_pmos ad=79.8f pd=0.8u as=0.1428p ps=1.52u w=0.42u l=0.13u
X476 a_58454_40850# vco_wob_0.vctl VSS VSS sg13_lv_nmos ad=65.99999f pd=0.74u as=0.102p ps=1.28u w=0.3u l=0.13u
X477 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.nQ a_62654_20215# VDD VDD sg13_lv_pmos ad=0.7616p pd=3.6u as=0.2163p ps=1.55u w=1.12u l=0.13u
X478 VDD a_62654_21971# a_62900_21935# VDD sg13_lv_pmos ad=0.2163p pd=1.55u as=79.8f ps=0.8u w=0.42u l=0.13u
X479 a_54504_22015# 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.D a_55086_21975# VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=50.4f ps=0.66u w=0.42u l=0.13u
X480 a_55770_40850# a_55831_40413# a_54489_40413# VSS sg13_lv_nmos ad=0.17p pd=1.68u as=0.11p ps=0.94u w=0.5u l=0.13u
X481 a_54602_21487# 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.Q 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.D VSS sg13_lv_nmos ad=88.8f pd=0.98u as=0.1628p ps=1.18u w=0.74u l=0.13u
X482 a_56039_25022# a_56013_24979# a_55941_24882# VSS sg13_lv_nmos ad=0.2307p pd=1.615u as=0.27427p ps=2.28u w=0.795u l=0.13u
X483 a_51685_23725# a_51648_24041# a_52119_23843# VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=47.25f ps=0.645u w=0.42u l=0.13u
X484 a_54898_22885# 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.Q a_54434_23148# VDD sg13_lv_pmos ad=0.1225p pd=1.245u as=0.34p ps=2.68u w=1u l=0.13u
X485 a_51693_23426# a_51631_22774# a_51684_22284# VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0.1428p ps=1.52u w=0.42u l=0.13u
X486 VSS a_56887_49467# VSS VSS sg13_lv_nmos ad=95f pd=0.88u as=0 ps=0 w=0.5u l=0.65u
X487 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.D a_61707_21488# a_61878_21130# VDD sg13_lv_pmos ad=0.3808p pd=2.92u as=0.2128p ps=1.5u w=1.12u l=0.13u
X488 VSS 3bit_freq_divider_1.dff_nclk_0.sg13g2_dfrbp_1_0.CLK a_64383_23628# VSS sg13_lv_nmos ad=0.1544p pd=1.235u as=0.2516p ps=2.16u w=0.74u l=0.13u
X489 VSS 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.Q a_53054_24999# VSS sg13_lv_nmos ad=0.15245p pd=1.17u as=88.8f ps=0.98u w=0.74u l=0.13u
X490 a_61887_20534# a_61691_20534# VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0.19p ps=1.38u w=1u l=0.13u
X491 VSS a_56887_49467# VSS VSS sg13_lv_nmos ad=95f pd=0.88u as=0 ps=0 w=0.5u l=0.65u
X492 VSS a_56887_49467# VSS VSS sg13_lv_nmos ad=95f pd=0.88u as=0 ps=0 w=0.5u l=0.65u
X493 a_64714_21300# 3bit_freq_divider_1.sg13g2_or3_1_0.A VDD VDD sg13_lv_pmos ad=0.22p pd=1.44u as=0.3822p ps=1.84u w=1u l=0.13u
X494 a_54504_20259# 3bit_freq_divider_0.dff_nclk_0.nCLK VDD VDD sg13_lv_pmos ad=79.8f pd=0.8u as=0.1428p ps=1.52u w=0.42u l=0.13u
X495 a_61707_21488# 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.Q a_61675_21130# VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0.1225p ps=1.245u w=1u l=0.13u
X496 VDD 3bit_freq_divider_1.dff_nclk_0.sg13g2_dfrbp_1_0.CLK a_64383_23628# VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0.34p ps=2.68u w=1u l=0.13u
X497 a_51684_22692# a_51631_22774# VSS VSS sg13_lv_nmos ad=0.2516p pd=2.16u as=0.1544p ps=1.235u w=0.74u l=0.13u
X498 a_57111_40283# a_53022_43738# VDD VDD sg13_lv_pmos ad=59.75f pd=0.745u as=59f ps=0.74u w=0.2u l=0.13u
X499 a_57112_40850# a_57173_40413# a_55831_40413# VSS sg13_lv_nmos ad=0.17p pd=1.68u as=0.11p ps=0.94u w=0.5u l=0.13u
X500 VDD a_53774_20178# a_53738_20514# VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0.34p ps=2.68u w=1u l=0.13u
X501 VDD a_51693_23075# a_51729_23026# VDD sg13_lv_pmos ad=0.11785p pd=1.025u as=51.45f ps=0.665u w=0.42u l=0.13u
X502 VSS charge_pump_0.vout VSS VSS sg13_lv_nmos ad=0.285p pd=1.88u as=0 ps=0 w=1.5u l=0.65u
X503 a_45451_28860# CLK_IN a_45579_29803# VSS sg13_lv_nmos ad=68.39999f pd=0.74u as=68.39999f ps=0.74u w=0.36u l=0.15u
X504 a_55345_21385# 3bit_freq_divider_0.freq_div_cell_0.Cout a_55485_21477# VSS sg13_lv_nmos ad=0.2176p pd=1.96u as=0.1216p ps=1.02u w=0.64u l=0.13u
X505 a_57173_40413# a_58515_40413# a_58454_40850# VSS sg13_lv_nmos ad=0.11p pd=0.94u as=0.17p ps=1.68u w=0.5u l=0.13u
X506 charge_pump_0.bias_p charge_pump_0.bias_n a_56742_53480# VSS sg13_lv_nmos ad=0.34p pd=2.68u as=0.34p ps=2.68u w=1u l=1u
X507 VSS a_56887_49467# VSS VSS sg13_lv_nmos ad=95f pd=0.88u as=0 ps=0 w=0.5u l=0.65u
X508 a_62270_22299# a_62119_22361# VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0.34p ps=2.68u w=1u l=0.13u
X509 VSS a_56887_49467# VSS VSS sg13_lv_nmos ad=95f pd=0.88u as=0 ps=0 w=0.5u l=0.65u
X510 a_64817_23685# a_64383_23434# a_64383_23889# VDD sg13_lv_pmos ad=43.05f pd=0.625u as=0.17695p ps=1.56u w=0.42u l=0.13u
X511 a_51648_24041# a_51631_22774# a_51693_23075# VDD sg13_lv_pmos ad=0.17695p pd=1.56u as=0.19p ps=1.38u w=1u l=0.13u
X512 VDD a_45658_27900# PFD_0.DOWN VDD sg13_lv_pmos ad=60.8f pd=0.7u as=0.1088p ps=1.32u w=0.32u l=0.15u
X513 3bit_freq_divider_1.freq_div_cell_0.Cout a_60967_23234# VDD VDD sg13_lv_pmos ad=0.3808p pd=2.92u as=0.1918p ps=1.5u w=1.12u l=0.13u
X514 a_64419_23844# 3bit_freq_divider_1.dff_nclk_0.nRST VSS VSS sg13_lv_nmos ad=47.25f pd=0.645u as=90.3f ps=0.85u w=0.42u l=0.13u
X515 3bit_freq_divider_1.sg13g2_or3_1_0.C Y0 a_63520_25000# VSS sg13_lv_nmos ad=0.1628p pd=1.18u as=88.8f ps=0.98u w=0.74u l=0.13u
X516 VSS a_64383_23889# a_64384_24445# VSS sg13_lv_nmos ad=0.14505p pd=1.15u as=0.187p ps=1.78u w=0.55u l=0.13u
X517 a_64384_21091# 3bit_freq_divider_1.sg13g2_or3_1_0.C a_64714_21414# VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0.1275p ps=1.255u w=1u l=0.13u
X518 VSS charge_pump_0.vout VSS VSS sg13_lv_nmos ad=0.285p pd=1.88u as=0 ps=0 w=1.5u l=0.65u
X519 VSS a_53968_20434# a_53899_20488# VSS sg13_lv_nmos ad=0.1825p pd=1.325u as=0.19397p ps=1.29u w=0.64u l=0.13u
X520 a_45451_28860# CLK_IN a_45579_29803# VSS sg13_lv_nmos ad=68.39999f pd=0.74u as=68.39999f ps=0.74u w=0.36u l=0.15u
X521 VDD 3bit_freq_divider_1.dff_nclk_0.nCLK a_61394_20220# VDD sg13_lv_pmos ad=0.1428p pd=1.52u as=79.8f ps=0.8u w=0.42u l=0.13u
X522 a_54489_40413# VSS cap_cmim l=6.99u w=6.99u
X523 VSS a_53065_23691# 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.nQ VSS sg13_lv_nmos ad=0.2516p pd=2.16u as=0.2775p ps=2.23u w=0.74u l=0.13u
X524 a_53899_20488# a_53774_20178# a_53065_20179# VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0.17695p ps=1.56u w=1u l=0.13u
X525 a_52074_23129# a_51693_23075# a_52074_23051# VSS sg13_lv_nmos ad=48.3f pd=0.65u as=54.6f ps=0.68u w=0.42u l=0.13u
X526 a_62324_23772# a_62270_24055# a_62246_23772# VSS sg13_lv_nmos ad=48.3f pd=0.65u as=54.6f ps=0.68u w=0.42u l=0.13u
X527 VDD CLK_IN a_45579_29803# VDD sg13_lv_pmos ad=60.8f pd=0.7u as=0.1088p ps=1.32u w=0.32u l=0.15u
X528 a_54352_24116# a_53899_24000# VDD VDD sg13_lv_pmos ad=51.45f pd=0.665u as=0.11785p ps=1.025u w=0.42u l=0.13u
X529 VDD X1 a_52924_22885# VDD sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X530 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.D 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.Q a_61972_21488# VSS sg13_lv_nmos ad=0.1628p pd=1.18u as=88.8f ps=0.98u w=0.74u l=0.13u
X531 VDD 3bit_freq_divider_1.freq_div_cell_0.Cin a_61878_22886# VDD sg13_lv_pmos ad=0.2128p pd=1.5u as=0.3808p ps=2.92u w=1.12u l=0.13u
X532 VSS a_53774_23690# a_53738_24026# VSS sg13_lv_nmos ad=0.1544p pd=1.235u as=0.2516p ps=2.16u w=0.74u l=0.13u
X533 a_54489_40413# a_55831_40413# a_55769_40283# VDD sg13_lv_pmos ad=0.11p pd=0.94u as=0.17p ps=1.68u w=0.5u l=0.13u
X534 a_61061_23234# 3bit_freq_divider_1.freq_div_cell_0.Cin a_60967_23234# VSS sg13_lv_nmos ad=0.1216p pd=1.02u as=0.2176p ps=1.96u w=0.64u l=0.13u
X535 a_55862_56737# charge_pump_0.bias_p charge_pump_0.bias_n VDD sg13_lv_pmos ad=0.38p pd=2.38u as=0.68p ps=4.68u w=2u l=1u
X536 a_62900_21935# a_62654_21971# a_63038_21971# VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=47.25f ps=0.645u w=0.42u l=0.13u
X537 a_63038_21971# 3bit_freq_divider_1.dff_nclk_0.nCLK VSS VSS sg13_lv_nmos ad=47.25f pd=0.645u as=90.3f ps=0.85u w=0.42u l=0.13u
X538 VSS charge_pump_0.vout VSS VSS sg13_lv_nmos ad=0.285p pd=1.88u as=0 ps=0 w=1.5u l=0.65u
X539 3bit_freq_divider_0.dff_nclk_0.D a_51648_24041# VSS VSS sg13_lv_nmos ad=0.2775p pd=2.23u as=0.2516p ps=2.16u w=0.74u l=0.13u
X540 a_51721_24988# a_51721_24988# a_52065_24890# VSS sg13_lv_nmos ad=0.102p pd=1.28u as=0.2307p ps=1.615u w=0.3u l=0.13u
X541 VSS a_55345_23141# 3bit_freq_divider_0.freq_div_cell_0.Cout VSS sg13_lv_nmos ad=0.1331p pd=1.12u as=0.2516p ps=2.16u w=0.74u l=0.13u
X542 a_52886_24904# X0 VSS VSS sg13_lv_nmos ad=0.17462p pd=1.185u as=0.15245p ps=1.17u w=0.55u l=0.13u
X543 VSS charge_pump_0.vout VSS VSS sg13_lv_nmos ad=0.285p pd=1.88u as=0 ps=0 w=1.5u l=0.65u
X544 a_55831_40413# a_57173_40413# a_57111_40283# VDD sg13_lv_pmos ad=0.11p pd=0.94u as=0.17p ps=1.68u w=0.5u l=0.13u
X545 a_54504_23771# 3bit_freq_divider_0.dff_nclk_0.nCLK VDD VDD sg13_lv_pmos ad=79.8f pd=0.8u as=0.1428p ps=1.52u w=0.42u l=0.13u
X546 a_62119_24117# a_61691_24046# a_61394_23732# VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0.1428p ps=1.52u w=0.42u l=0.13u
X547 VSS 3bit_freq_divider_1.dff_nclk_0.nCLK a_61488_23732# VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=50.4f ps=0.66u w=0.42u l=0.13u
X548 3bit_freq_divider_0.EN nEN VSS VSS sg13_lv_nmos ad=0.259p pd=2.18u as=0.259p ps=2.18u w=0.74u l=0.13u
X549 VSS charge_pump_0.vout VSS VSS sg13_lv_nmos ad=0.285p pd=1.88u as=0 ps=0 w=1.5u l=0.65u
X550 a_59799_40285# a_53022_43738# VDD VDD sg13_lv_pmos ad=59.75f pd=0.745u as=59f ps=0.74u w=0.2u l=0.13u
X551 a_53899_20488# a_53738_20514# a_53065_20179# VSS sg13_lv_nmos ad=0.19397p pd=1.29u as=0.2017p ps=1.48u w=0.64u l=0.13u
X552 VSS PFD_0.VCO_CLK a_45451_28860# VSS sg13_lv_nmos ad=0.1224p pd=1.4u as=0.1224p ps=1.4u w=0.36u l=0.15u
X553 VSS a_46817_27899# a_45658_27900# VSS sg13_lv_nmos ad=0.1224p pd=1.4u as=0.1224p ps=1.4u w=0.36u l=0.15u
X554 a_53054_21487# X2 3bit_freq_divider_0.sg13g2_or3_1_0.A VSS sg13_lv_nmos ad=88.8f pd=0.98u as=0.1628p ps=1.18u w=0.74u l=0.13u
X555 a_53350_22885# X1 a_52886_23148# VDD sg13_lv_pmos ad=0.1225p pd=1.245u as=0.34p ps=2.68u w=1u l=0.13u
X556 VSS vco_wob_0.vctl a_57311_42591# VSS sg13_lv_nmos ad=0.102p pd=1.28u as=65.99999f ps=0.74u w=0.3u l=0.13u
X557 a_62900_23691# 3bit_freq_divider_1.dff_nclk_0.nCLK VDD VDD sg13_lv_pmos ad=79.8f pd=0.8u as=79.8f ps=0.8u w=0.42u l=0.13u
X558 a_53774_23690# 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.sg13g2_dfrbp_1_0.CLK VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0.19p ps=1.38u w=1u l=0.13u
X559 a_57311_42591# a_55836_43159# a_57178_43159# VSS sg13_lv_nmos ad=0.17p pd=1.68u as=0.11p ps=0.94u w=0.5u l=0.13u
X560 a_58653_42591# vco_wob_0.vctl VSS VSS sg13_lv_nmos ad=65.99999f pd=0.74u as=0.102p ps=1.28u w=0.3u l=0.13u
X561 a_55831_40413# a_57173_40413# a_57111_40283# VDD sg13_lv_pmos ad=0.1106p pd=0.945u as=0.11p ps=0.94u w=0.5u l=0.13u
X562 a_60967_21478# 3bit_freq_divider_1.freq_div_cell_0.Cout VDD VDD sg13_lv_pmos ad=0.1596p pd=1.22u as=0.2856p ps=2.36u w=0.84u l=0.13u
X563 VSS a_62900_21935# a_62848_21971# VSS sg13_lv_nmos ad=90.3f pd=0.85u as=54.6f ps=0.68u w=0.42u l=0.13u
X564 a_58426_43159# a_57178_43159# 3bit_freq_divider_0.CLK_IN VDD sg13_lv_pmos ad=0.17p pd=1.68u as=0.11p ps=0.94u w=0.5u l=0.13u
X565 3bit_freq_divider_0.CLK_IN a_57178_43159# a_58653_42591# VSS sg13_lv_nmos ad=0.11p pd=0.94u as=0.17p ps=1.68u w=0.5u l=0.13u
X566 VDD 3bit_freq_divider_0.dff_nclk_0.nCLK a_53968_20434# VDD sg13_lv_pmos ad=0.11785p pd=1.025u as=0.1533p ps=1.57u w=0.42u l=0.13u
X567 a_62119_24117# a_61887_24046# a_61394_23732# VDD sg13_lv_pmos ad=79.8f pd=0.8u as=0.1428p ps=1.52u w=0.42u l=0.13u
X568 a_54747_49259# charge_pump_0.bias_n VSS VSS sg13_lv_nmos ad=0.207p pd=1.545u as=0.408p ps=3.08u w=1.2u l=0.13u
X569 VDD a_53022_43738# a_54400_43159# VDD sg13_lv_pmos ad=59f pd=0.74u as=59.75f ps=0.745u w=0.2u l=0.13u
X570 VDD a_53022_43738# a_53022_43738# VDD sg13_lv_pmos ad=59f pd=0.74u as=59f ps=0.74u w=0.2u l=0.13u
X571 VSS 3bit_freq_divider_1.dff_nclk_0.nCLK a_62324_20260# VSS sg13_lv_nmos ad=0.1825p pd=1.325u as=48.3f ps=0.65u w=0.42u l=0.13u
X572 a_62848_21971# a_61691_22290# a_62654_21971# VSS sg13_lv_nmos ad=54.6f pd=0.68u as=0.2017p ps=1.48u w=0.42u l=0.13u
X573 a_63255_23244# Y1 a_63223_22886# VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0.1225p ps=1.245u w=1u l=0.13u
X574 a_53774_23690# 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.sg13g2_dfrbp_1_0.CLK VSS VSS sg13_lv_nmos ad=0.2516p pd=2.16u as=0.1544p ps=1.235u w=0.74u l=0.13u
X575 VSS 3bit_freq_divider_0.sg13g2_tiehi_1.L_HI a_54434_24904# VSS sg13_lv_nmos ad=0.374p pd=2.46u as=0.17462p ps=1.185u w=0.55u l=0.13u
X576 a_60385_24558# a_60385_24947# a_60385_24717# VDD sg13_lv_pmos ad=0.4657p pd=2.54u as=0.2442p ps=2.06u w=0.66u l=0.13u
X577 VSS Y1 a_63255_23244# VSS sg13_lv_nmos ad=0.15245p pd=1.17u as=0.17462p ps=1.185u w=0.55u l=0.13u
X578 a_58453_40283# a_58515_40413# a_57173_40413# VDD sg13_lv_pmos ad=0.17p pd=1.68u as=0.1106p ps=0.945u w=0.5u l=0.13u
X579 a_46749_30782# CLK_IN CLK_IN VDD sg13_lv_pmos ad=0.1088p pd=1.32u as=60.8f ps=0.7u w=0.32u l=0.15u
X580 a_61675_21130# 3bit_freq_divider_1.freq_div_cell_0.Cout VDD VDD sg13_lv_pmos ad=0.1225p pd=1.245u as=0.36p ps=2.72u w=1u l=0.13u
X581 a_52119_23653# a_51631_22774# a_51648_24041# VSS sg13_lv_nmos ad=54.6f pd=0.68u as=0.2017p ps=1.48u w=0.42u l=0.13u
X582 a_52950_22157# a_53065_21935# VDD VDD sg13_lv_pmos ad=0.2856p pd=2.36u as=0.2016p ps=1.5u w=0.84u l=0.13u
X583 PFD_0.VCO_CLK a_51648_24438# VDD VDD sg13_lv_pmos ad=0.3808p pd=2.92u as=0.2016p ps=1.5u w=1.12u l=0.13u
X584 3bit_freq_divider_1.dff_nclk_0.D a_64383_23889# VSS VSS sg13_lv_nmos ad=0.2775p pd=2.23u as=0.2516p ps=2.16u w=0.74u l=0.13u
X585 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 3bit_freq_divider_1.sg13g2_nand2_1_0.Y VDD VDD sg13_lv_pmos ad=0.392p pd=2.94u as=0.392p ps=2.94u w=1.12u l=0.13u
X586 VDD a_62900_20179# a_62879_20613# VDD sg13_lv_pmos ad=79.8f pd=0.8u as=43.05f ps=0.625u w=0.42u l=0.13u
X587 a_55345_21385# 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.Q VDD VDD sg13_lv_pmos ad=0.1596p pd=1.22u as=0.1918p ps=1.5u w=0.84u l=0.13u
X588 VDD a_53065_20179# 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.nQ VDD sg13_lv_pmos ad=0.2163p pd=1.55u as=0.7616p ps=3.6u w=1.12u l=0.13u
X589 a_51648_21103# 3bit_freq_divider_0.sg13g2_or3_1_0.A VSS VSS sg13_lv_nmos ad=0.198p pd=1.27u as=0.13395p ps=1.12u w=0.55u l=0.13u
X590 VSS a_51648_21103# 3bit_freq_divider_0.dff_nclk_0.nCLK VSS sg13_lv_nmos ad=0.13395p pd=1.12u as=0.2516p ps=2.16u w=0.74u l=0.13u
X591 a_52944_43077# a_53147_40413# a_53085_40283# VDD sg13_lv_pmos ad=0.1106p pd=0.945u as=0.11p ps=0.94u w=0.5u l=0.13u
X592 a_59799_40285# 3bit_freq_divider_0.CLK_IN a_58515_40413# VDD sg13_lv_pmos ad=0.11p pd=0.94u as=0.11p ps=0.94u w=0.5u l=0.13u
X593 a_53065_23691# a_53738_24026# a_53702_24124# VDD sg13_lv_pmos ad=0.17695p pd=1.56u as=43.05f ps=0.625u w=0.42u l=0.13u
X594 a_54504_22015# a_53738_22270# a_53968_22190# VDD sg13_lv_pmos ad=0.1428p pd=1.52u as=79.8f ps=0.8u w=0.42u l=0.13u
X595 VDD a_53022_43738# a_54400_43159# VDD sg13_lv_pmos ad=0.104p pd=1.34u as=59f ps=0.74u w=0.2u l=0.13u
X596 VDD a_62654_21971# a_63463_21972# VDD sg13_lv_pmos ad=0.2016p pd=1.5u as=0.2856p ps=2.36u w=0.84u l=0.13u
X597 a_47954_28913# PFD_0.VCO_CLK VDD VDD sg13_lv_pmos ad=0.1088p pd=1.32u as=60.8f ps=0.7u w=0.32u l=0.15u
X598 VDD 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.Q a_60967_24990# VDD sg13_lv_pmos ad=0.1918p pd=1.5u as=0.1596p ps=1.22u w=0.84u l=0.13u
X599 a_52950_20401# a_53065_20179# VSS VSS sg13_lv_nmos ad=0.187p pd=1.78u as=0.14505p ps=1.15u w=0.55u l=0.13u
X600 a_53086_40850# vco_wob_0.vctl VSS VSS sg13_lv_nmos ad=65.99999f pd=0.74u as=0.102p ps=1.28u w=0.3u l=0.13u
X601 a_62246_23772# a_61887_24046# a_62119_24117# VSS sg13_lv_nmos ad=54.6f pd=0.68u as=79.8f ps=0.8u w=0.42u l=0.13u
X602 VDD 3bit_freq_divider_0.freq_div_cell_0.Cin a_54898_22885# VDD sg13_lv_pmos ad=0.36p pd=2.72u as=0.1225p ps=1.245u w=1u l=0.13u
X603 VDD a_53022_43738# a_57111_40283# VDD sg13_lv_pmos ad=0.104p pd=1.34u as=59.75f ps=0.745u w=0.2u l=0.13u
X604 a_48909_28913# PFD_0.VCO_CLK a_47954_28913# VSS sg13_lv_nmos ad=68.39999f pd=0.74u as=68.39999f ps=0.74u w=0.36u l=0.15u
X605 VSS 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.Q a_52886_21392# VSS sg13_lv_nmos ad=0.374p pd=2.46u as=0.17462p ps=1.185u w=0.55u l=0.13u
X606 a_55345_24897# 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.Q VDD VDD sg13_lv_pmos ad=0.1596p pd=1.22u as=0.1918p ps=1.5u w=0.84u l=0.13u
X607 VSS charge_pump_0.vout VSS VSS sg13_lv_nmos ad=0.285p pd=1.88u as=0 ps=0 w=1.5u l=0.65u
X608 a_58453_40283# a_53022_43738# VDD VDD sg13_lv_pmos ad=59.75f pd=0.745u as=59f ps=0.74u w=0.2u l=0.13u
X609 3bit_freq_divider_0.sg13g2_or3_1_0.B a_52886_23148# VSS VSS sg13_lv_nmos ad=0.1628p pd=1.18u as=0.3108p ps=2.32u w=0.74u l=0.13u
X610 VSS a_62654_20215# a_63463_20216# VSS sg13_lv_nmos ad=0.14505p pd=1.15u as=0.187p ps=1.78u w=0.55u l=0.13u
X611 a_63255_21488# 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.Q VSS VSS sg13_lv_nmos ad=0.17462p pd=1.185u as=0.374p ps=2.46u w=0.55u l=0.13u
X612 a_54252_22015# 3bit_freq_divider_0.dff_nclk_0.nCLK VSS VSS sg13_lv_nmos ad=48.3f pd=0.65u as=0.1825p ps=1.325u w=0.42u l=0.13u
X613 a_63426_22886# Y1 VDD VDD sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X614 VDD a_53022_43738# a_55742_43159# VDD sg13_lv_pmos ad=0.104p pd=1.34u as=59f ps=0.74u w=0.2u l=0.13u
X615 a_51685_23725# 3bit_freq_divider_0.dff_nclk_0.nRST VDD VDD sg13_lv_pmos ad=79.8f pd=0.8u as=79.8f ps=0.8u w=0.42u l=0.13u
X616 a_53539_20214# a_53065_20179# a_53445_20214# VSS sg13_lv_nmos ad=47.25f pd=0.645u as=0.1428p ps=1.52u w=0.42u l=0.13u
X617 VSS 3bit_freq_divider_0.dff_nclk_0.nCLK a_53539_20214# VSS sg13_lv_nmos ad=90.3f pd=0.85u as=47.25f ps=0.645u w=0.42u l=0.13u
X618 VDD 3bit_freq_divider_0.EN 3bit_freq_divider_0.sg13g2_nand2_1_0.Y VDD sg13_lv_pmos ad=0.3808p pd=2.92u as=0.2128p ps=1.5u w=1.12u l=0.13u
X619 a_54504_22015# a_53774_21934# a_53968_22190# VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=79.8f ps=0.8u w=0.42u l=0.13u
X620 3bit_freq_divider_1.sg13g2_or3_1_0.A a_63255_21488# a_63426_21130# VDD sg13_lv_pmos ad=0.3808p pd=2.92u as=0.2128p ps=1.5u w=1.12u l=0.13u
X621 a_52924_21129# a_52886_21392# 3bit_freq_divider_0.sg13g2_or3_1_0.A VDD sg13_lv_pmos ad=0.2128p pd=1.5u as=0.3808p ps=2.92u w=1.12u l=0.13u
X622 VDD 3bit_freq_divider_1.dff_nclk_0.nCLK a_61394_21976# VDD sg13_lv_pmos ad=0.1428p pd=1.52u as=79.8f ps=0.8u w=0.42u l=0.13u
X623 a_57178_43159# a_55836_43159# a_57084_43159# VDD sg13_lv_pmos ad=0.11p pd=0.94u as=0.11p ps=0.94u w=0.5u l=0.13u
X624 VSS 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.sg13g2_dfrbp_1_0.CLK a_61691_20534# VSS sg13_lv_nmos ad=0.1544p pd=1.235u as=0.2516p ps=2.16u w=0.74u l=0.13u
X625 a_53968_20434# a_53774_20178# a_54352_20604# VDD sg13_lv_pmos ad=79.8f pd=0.8u as=51.45f ps=0.665u w=0.42u l=0.13u
X626 a_64419_23326# a_64383_23300# VSS VSS sg13_lv_nmos ad=0.19397p pd=1.29u as=0.1825p ps=1.325u w=0.64u l=0.13u
X627 a_52944_43077# a_53147_40413# a_53086_40850# VSS sg13_lv_nmos ad=0.11p pd=0.94u as=0.17p ps=1.68u w=0.5u l=0.13u
X628 3bit_freq_divider_1.sg13g2_nand2_1_0.Y 3bit_freq_divider_0.EN VDD VDD sg13_lv_pmos ad=0.2128p pd=1.5u as=0.3808p ps=2.92u w=1.12u l=0.13u
X629 VSS charge_pump_0.vout VSS VSS sg13_lv_nmos ad=0.285p pd=1.88u as=0 ps=0 w=1.5u l=0.65u
X630 a_47954_28913# PFD_0.VCO_CLK a_46817_27899# VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0.1428p ps=1.52u w=0.42u l=0.15u
X631 a_62270_22299# a_62119_22361# VSS VSS sg13_lv_nmos ad=0.19397p pd=1.29u as=0.1825p ps=1.325u w=0.64u l=0.13u
X632 a_62900_23691# a_62654_23727# a_63038_23727# VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=47.25f ps=0.645u w=0.42u l=0.13u
X633 a_63038_23727# 3bit_freq_divider_1.dff_nclk_0.nCLK VSS VSS sg13_lv_nmos ad=47.25f pd=0.645u as=90.3f ps=0.85u w=0.42u l=0.13u
X634 VDD a_53022_43738# a_53022_43738# VDD sg13_lv_pmos ad=0.104p pd=1.34u as=59.75f ps=0.745u w=0.2u l=0.13u
X635 a_52924_24641# a_52886_24904# 3bit_freq_divider_0.sg13g2_or3_1_0.C VDD sg13_lv_pmos ad=0.2128p pd=1.5u as=0.3808p ps=2.92u w=1.12u l=0.13u
X636 a_56137_24678# a_56137_24678# a_56039_25022# VSS sg13_lv_nmos ad=0.102p pd=1.28u as=0.2307p ps=1.615u w=0.3u l=0.13u
X637 a_45579_29803# CLK_IN a_45451_28860# VSS sg13_lv_nmos ad=68.39999f pd=0.74u as=0.1224p ps=1.4u w=0.36u l=0.15u
X638 VSS a_45658_27900# PFD_0.DOWN VSS sg13_lv_nmos ad=0.1632p pd=1.64u as=0.1632p ps=1.64u w=0.48u l=0.15u
X639 a_52944_43077# VSS cap_cmim l=6.99u w=6.99u
X640 a_53702_22368# a_53445_21970# VDD VDD sg13_lv_pmos ad=43.05f pd=0.625u as=79.8f ps=0.8u w=0.42u l=0.13u
X641 a_63520_23244# 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.Q VSS VSS sg13_lv_nmos ad=88.8f pd=0.98u as=0.15245p ps=1.17u w=0.74u l=0.13u
X642 a_61707_23244# 3bit_freq_divider_1.freq_div_cell_0.Cin VSS VSS sg13_lv_nmos ad=0.17462p pd=1.185u as=0.374p ps=2.46u w=0.55u l=0.13u
X643 a_51759_25014# a_51721_24988# a_51600_24907# VDD sg13_lv_pmos ad=0.2442p pd=2.06u as=0.4657p ps=2.54u w=0.66u l=0.13u
X644 VDD a_53968_23946# a_53899_24000# VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0.19p ps=1.38u w=1u l=0.13u
X645 VDD 3bit_freq_divider_0.freq_div_cell_0.Cout a_55345_21385# VDD sg13_lv_pmos ad=0.2856p pd=2.36u as=0.1596p ps=1.22u w=0.84u l=0.13u
X646 VSS 3bit_freq_divider_0.freq_div_cell_0.Cout a_54602_21487# VSS sg13_lv_nmos ad=0.15245p pd=1.17u as=88.8f ps=0.98u w=0.74u l=0.13u
X647 VSS a_56887_49467# VSS VSS sg13_lv_nmos ad=95f pd=0.88u as=0 ps=0 w=0.5u l=0.65u
X648 a_53058_43159# a_53022_43738# VDD VDD sg13_lv_pmos ad=59f pd=0.74u as=59f ps=0.74u w=0.2u l=0.13u
X649 VSS a_64384_21091# 3bit_freq_divider_1.dff_nclk_0.nCLK VSS sg13_lv_nmos ad=0.13395p pd=1.12u as=0.2516p ps=2.16u w=0.74u l=0.13u
X650 VDD a_62270_22299# a_62221_22361# VDD sg13_lv_pmos ad=0.11785p pd=1.025u as=51.45f ps=0.665u w=0.42u l=0.13u
X651 VSS vco_wob_0.vctl a_54627_42591# VSS sg13_lv_nmos ad=0.102p pd=1.28u as=65.99999f ps=0.74u w=0.3u l=0.13u
X652 a_51721_23684# a_51684_22692# a_51648_24041# VDD sg13_lv_pmos ad=43.05f pd=0.625u as=0.17695p ps=1.56u w=0.42u l=0.13u
X653 a_54627_42591# a_53152_43159# a_54494_43159# VSS sg13_lv_nmos ad=0.17p pd=1.68u as=0.11p ps=0.94u w=0.5u l=0.13u
X654 a_51684_22284# 3bit_freq_divider_0.dff_nclk_0.D VDD VDD sg13_lv_pmos ad=79.8f pd=0.8u as=0.1428p ps=1.52u w=0.42u l=0.13u
X655 a_61887_24046# a_61691_24046# VSS VSS sg13_lv_nmos ad=0.2516p pd=2.16u as=0.1544p ps=1.235u w=0.74u l=0.13u
X656 VDD a_53065_23691# 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.nQ VDD sg13_lv_pmos ad=0.2163p pd=1.55u as=0.7616p ps=3.6u w=1.12u l=0.13u
X657 a_53445_20214# a_53065_20179# VDD VDD sg13_lv_pmos ad=79.8f pd=0.8u as=0.2163p ps=1.55u w=0.42u l=0.13u
X658 VSS a_56887_49467# VSS VSS sg13_lv_nmos ad=95f pd=0.88u as=0 ps=0 w=0.5u l=0.65u
X659 VDD 3bit_freq_divider_0.sg13g2_tiehi_1.L_HI a_55345_24897# VDD sg13_lv_pmos ad=0.2856p pd=2.36u as=0.1596p ps=1.22u w=0.84u l=0.13u
X660 3bit_freq_divider_1.sg13g2_or3_1_0.A Y2 a_63520_21488# VSS sg13_lv_nmos ad=0.1628p pd=1.18u as=88.8f ps=0.98u w=0.74u l=0.13u
X661 VDD 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.Q a_54472_22885# VDD sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X662 CLK_OUT a_64384_24445# VDD VDD sg13_lv_pmos ad=0.3808p pd=2.92u as=0.2016p ps=1.5u w=1.12u l=0.13u
X663 VSS a_56887_49467# VSS VSS sg13_lv_nmos ad=95f pd=0.88u as=0 ps=0 w=0.5u l=0.65u
X664 a_53065_20179# a_53774_20178# a_53722_20214# VSS sg13_lv_nmos ad=0.2017p pd=1.48u as=54.6f ps=0.68u w=0.42u l=0.13u
X665 a_64424_22200# 3bit_freq_divider_1.dff_nclk_0.D VDD VDD sg13_lv_pmos ad=79.8f pd=0.8u as=0.1428p ps=1.52u w=0.42u l=0.13u
X666 a_63223_22886# 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.Q VDD VDD sg13_lv_pmos ad=0.1225p pd=1.245u as=0.36p ps=2.72u w=1u l=0.13u
X667 a_61488_21976# 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.D a_61394_21976# VSS sg13_lv_nmos ad=50.4f pd=0.66u as=0.1428p ps=1.52u w=0.42u l=0.13u
X668 VSS a_62900_23691# a_62848_23727# VSS sg13_lv_nmos ad=90.3f pd=0.85u as=54.6f ps=0.68u w=0.42u l=0.13u
X669 a_53722_20214# a_53445_20214# VSS VSS sg13_lv_nmos ad=54.6f pd=0.68u as=90.3f ps=0.85u w=0.42u l=0.13u
X670 a_64383_23706# a_64383_23889# a_64419_23844# VSS sg13_lv_nmos ad=0.1428p pd=1.52u as=47.25f ps=0.645u w=0.42u l=0.13u
X671 VSS 3bit_freq_divider_1.dff_nclk_0.nCLK a_62324_22016# VSS sg13_lv_nmos ad=0.1825p pd=1.325u as=48.3f ps=0.65u w=0.42u l=0.13u
X672 a_62848_23727# a_61691_24046# a_62654_23727# VSS sg13_lv_nmos ad=54.6f pd=0.68u as=0.2017p ps=1.48u w=0.42u l=0.13u
X673 VDD charge_pump_0.bias_p a_54842_49733# VDD sg13_lv_pmos ad=0.1005p pd=1.34u as=55.5f ps=0.74u w=0.15u l=0.13u
X674 VSS a_56887_49467# VSS VSS sg13_lv_nmos ad=95f pd=0.88u as=0 ps=0 w=0.5u l=0.65u
X675 a_46817_27899# PFD_0.VCO_CLK PFD_0.VCO_CLK VDD sg13_lv_pmos ad=0.1088p pd=1.32u as=60.8f ps=0.7u w=0.32u l=0.15u
X676 a_57173_40413# a_58515_40413# a_58453_40283# VDD sg13_lv_pmos ad=0.1106p pd=0.945u as=0.11p ps=0.94u w=0.5u l=0.13u
X677 a_64384_21091# 3bit_freq_divider_1.sg13g2_or3_1_0.C VSS VSS sg13_lv_nmos ad=0.187p pd=1.78u as=0.1045p ps=0.93u w=0.55u l=0.13u
X678 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 3bit_freq_divider_1.sg13g2_nand2_1_0.Y VSS VSS sg13_lv_nmos ad=0.259p pd=2.18u as=0.259p ps=2.18u w=0.74u l=0.13u
X679 VSS charge_pump_0.vout VSS VSS sg13_lv_nmos ad=0.51p pd=3.68u as=0 ps=0 w=1.5u l=0.65u
X680 a_53285_42591# vco_wob_0.vctl VSS VSS sg13_lv_nmos ad=65.99999f pd=0.74u as=0.102p ps=1.28u w=0.3u l=0.13u
X681 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.D a_54434_24904# VSS VSS sg13_lv_nmos ad=0.1628p pd=1.18u as=0.3108p ps=2.32u w=0.74u l=0.13u
X682 a_54504_23771# a_53738_24026# a_53968_23946# VDD sg13_lv_pmos ad=0.1428p pd=1.52u as=79.8f ps=0.8u w=0.42u l=0.13u
X683 a_61878_22886# 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.Q VDD VDD sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2128p ps=1.5u w=1.12u l=0.13u
X684 CLK_IN CLK_IN a_46749_30782# VDD sg13_lv_pmos ad=60.8f pd=0.7u as=0.1088p ps=1.32u w=0.32u l=0.15u
X685 a_53058_43159# a_52944_43077# a_53152_43159# VDD sg13_lv_pmos ad=0.17p pd=1.68u as=0.11p ps=0.94u w=0.5u l=0.13u
X686 a_53152_43159# a_52944_43077# a_53285_42591# VSS sg13_lv_nmos ad=0.11p pd=0.94u as=0.17p ps=1.68u w=0.5u l=0.13u
X687 a_54434_21392# 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.Q VSS VSS sg13_lv_nmos ad=0.17462p pd=1.185u as=0.15245p ps=1.17u w=0.55u l=0.13u
X688 VSS a_63255_25000# 3bit_freq_divider_1.sg13g2_or3_1_0.C VSS sg13_lv_nmos ad=0.3108p pd=2.32u as=0.1628p ps=1.18u w=0.74u l=0.13u
X689 a_47954_28913# PFD_0.VCO_CLK a_48909_28913# VSS sg13_lv_nmos ad=68.39999f pd=0.74u as=68.39999f ps=0.74u w=0.36u l=0.15u
X690 VDD 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.Q a_63426_24642# VDD sg13_lv_pmos ad=0.2128p pd=1.5u as=0.3808p ps=2.92u w=1.12u l=0.13u
X691 3bit_freq_divider_1.freq_div_cell_1.Cout a_60967_21478# VSS VSS sg13_lv_nmos ad=0.2516p pd=2.16u as=0.1331p ps=1.12u w=0.74u l=0.13u
X692 a_53085_40283# a_53147_40413# a_52944_43077# VDD sg13_lv_pmos ad=0.17p pd=1.68u as=0.1106p ps=0.945u w=0.5u l=0.13u
X693 a_54472_22885# 3bit_freq_divider_0.freq_div_cell_0.Cin VDD VDD sg13_lv_pmos ad=0.3808p pd=2.92u as=0.2128p ps=1.5u w=1.12u l=0.13u
X694 VSS charge_pump_0.vout VSS VSS sg13_lv_nmos ad=0.285p pd=1.88u as=0 ps=0 w=1.5u l=0.65u
X695 a_64383_23300# 3bit_freq_divider_1.dff_nclk_0.nRST VDD VDD sg13_lv_pmos ad=0.1533p pd=1.57u as=0.11785p ps=1.025u w=0.42u l=0.13u
X696 a_55769_40283# a_55831_40413# a_54489_40413# VDD sg13_lv_pmos ad=0.11p pd=0.94u as=0.11p ps=0.94u w=0.5u l=0.13u
X697 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.Q a_63463_21972# VSS VSS sg13_lv_nmos ad=0.2516p pd=2.16u as=0.14505p ps=1.15u w=0.74u l=0.13u
X698 a_54428_40850# vco_wob_0.vctl VSS VSS sg13_lv_nmos ad=65.99999f pd=0.74u as=0.102p ps=1.28u w=0.3u l=0.13u
X699 VDD PFD_0.VCO_CLK a_47954_28913# VDD sg13_lv_pmos ad=60.8f pd=0.7u as=0.1088p ps=1.32u w=0.32u l=0.15u
X700 a_54352_20604# a_53899_20488# VDD VDD sg13_lv_pmos ad=51.45f pd=0.665u as=0.11785p ps=1.025u w=0.42u l=0.13u
X701 charge_pump_0.vout a_56887_49467# rhigh l=0.96u w=0.5u
X702 a_55836_43159# a_54494_43159# a_55742_43159# VDD sg13_lv_pmos ad=0.11p pd=0.94u as=0.11p ps=0.94u w=0.5u l=0.13u
X703 VDD a_53022_43738# a_58453_40283# VDD sg13_lv_pmos ad=0.104p pd=1.34u as=59.75f ps=0.745u w=0.2u l=0.13u
X704 3bit_freq_divider_1.freq_div_cell_0.Cin a_60967_24990# VSS VSS sg13_lv_nmos ad=0.2516p pd=2.16u as=0.1331p ps=1.12u w=0.74u l=0.13u
X705 VSS 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.Q a_53054_21487# VSS sg13_lv_nmos ad=0.15245p pd=1.17u as=88.8f ps=0.98u w=0.74u l=0.13u
X706 VSS 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK a_61691_22290# VSS sg13_lv_nmos ad=0.1544p pd=1.235u as=0.2516p ps=2.16u w=0.74u l=0.13u
X707 VDD 3bit_freq_divider_0.dff_nclk_0.nCLK a_53445_23726# VDD sg13_lv_pmos ad=79.8f pd=0.8u as=79.8f ps=0.8u w=0.42u l=0.13u
X708 VSS charge_pump_0.vout VSS VSS sg13_lv_nmos ad=0.285p pd=1.88u as=0 ps=0 w=1.5u l=0.65u
X709 a_54472_21129# a_54434_21392# 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.D VDD sg13_lv_pmos ad=0.2128p pd=1.5u as=0.3808p ps=2.92u w=1.12u l=0.13u
X710 VDD 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.Q a_53350_21129# VDD sg13_lv_pmos ad=0.36p pd=2.72u as=0.1225p ps=1.245u w=1u l=0.13u
X711 a_57111_40283# a_57173_40413# a_55831_40413# VDD sg13_lv_pmos ad=0.11p pd=0.94u as=0.11p ps=0.94u w=0.5u l=0.13u
X712 a_52065_24890# a_51759_25014# a_51622_24863# VSS sg13_lv_nmos ad=0.2307p pd=1.615u as=0.27427p ps=2.28u w=0.795u l=0.13u
X713 a_62270_24055# a_62119_24117# VSS VSS sg13_lv_nmos ad=0.19397p pd=1.29u as=0.1825p ps=1.325u w=0.64u l=0.13u
X714 a_58426_43159# a_53022_43738# VDD VDD sg13_lv_pmos ad=59f pd=0.74u as=59f ps=0.74u w=0.2u l=0.13u
X715 a_57173_40413# a_58515_40413# a_58453_40283# VDD sg13_lv_pmos ad=0.11p pd=0.94u as=0.17p ps=1.68u w=0.5u l=0.13u
X716 VDD a_53022_43738# a_59799_40285# VDD sg13_lv_pmos ad=59f pd=0.74u as=59f ps=0.74u w=0.2u l=0.13u
X717 a_64383_23889# a_64383_23434# a_64419_23326# VSS sg13_lv_nmos ad=0.2017p pd=1.48u as=0.19397p ps=1.29u w=0.64u l=0.13u
X718 a_53085_40283# a_53022_43738# VDD VDD sg13_lv_pmos ad=59.75f pd=0.745u as=59f ps=0.74u w=0.2u l=0.13u
X719 VDD a_53022_43738# a_54427_40283# VDD sg13_lv_pmos ad=59f pd=0.74u as=59f ps=0.74u w=0.2u l=0.13u
X720 VDD a_53022_43738# a_59799_40285# VDD sg13_lv_pmos ad=0.104p pd=1.34u as=59.75f ps=0.745u w=0.2u l=0.13u
X721 a_62221_22361# a_61691_22290# a_62119_22361# VDD sg13_lv_pmos ad=51.45f pd=0.665u as=79.8f ps=0.8u w=0.42u l=0.13u
X722 a_56742_53480# VSS rhigh l=12u w=1u
X723 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.Q a_63463_23728# VDD VDD sg13_lv_pmos ad=0.3808p pd=2.92u as=0.2016p ps=1.5u w=1.12u l=0.13u
X724 a_53147_40413# a_54489_40413# a_54428_40850# VSS sg13_lv_nmos ad=0.11p pd=0.94u as=0.17p ps=1.68u w=0.5u l=0.13u
X725 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.D a_61707_23244# a_61878_22886# VDD sg13_lv_pmos ad=0.3808p pd=2.92u as=0.2128p ps=1.5u w=1.12u l=0.13u
X726 VDD a_62270_24055# a_62221_24117# VDD sg13_lv_pmos ad=0.11785p pd=1.025u as=51.45f ps=0.665u w=0.42u l=0.13u
X727 VSS charge_pump_0.vout VSS VSS sg13_lv_nmos ad=0.285p pd=1.88u as=0 ps=0 w=1.5u l=0.65u
X728 a_54472_24641# a_54434_24904# 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.D VDD sg13_lv_pmos ad=0.2128p pd=1.5u as=0.3808p ps=2.92u w=1.12u l=0.13u
X729 VDD 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.Q a_53350_24641# VDD sg13_lv_pmos ad=0.36p pd=2.72u as=0.1225p ps=1.245u w=1u l=0.13u
X730 a_53058_43159# a_52944_43077# a_53152_43159# VDD sg13_lv_pmos ad=0.11p pd=0.94u as=0.1106p ps=0.945u w=0.5u l=0.13u
X731 VDD 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.D a_54504_20259# VDD sg13_lv_pmos ad=0.1428p pd=1.52u as=79.8f ps=0.8u w=0.42u l=0.13u
X732 a_61707_23244# 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.Q a_61675_22886# VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0.1225p ps=1.245u w=1u l=0.13u
X733 a_64419_23326# a_64383_23300# VDD VDD sg13_lv_pmos ad=0.19p pd=1.38u as=0.34p ps=2.68u w=1u l=0.13u
X734 a_51708_21413# 3bit_freq_divider_0.sg13g2_or3_1_0.B a_51708_21299# VDD sg13_lv_pmos ad=0.1275p pd=1.255u as=0.22p ps=1.44u w=1u l=0.13u
X735 VSS 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.Q a_61707_23244# VSS sg13_lv_nmos ad=0.15245p pd=1.17u as=0.17462p ps=1.185u w=0.55u l=0.13u
X736 VSS a_53065_20179# 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.nQ VSS sg13_lv_nmos ad=0.2516p pd=2.16u as=0.2775p ps=2.23u w=0.74u l=0.13u
X737 a_62324_20260# a_62270_20543# a_62246_20260# VSS sg13_lv_nmos ad=48.3f pd=0.65u as=54.6f ps=0.68u w=0.42u l=0.13u
X738 a_62900_20179# 3bit_freq_divider_1.dff_nclk_0.nCLK VDD VDD sg13_lv_pmos ad=79.8f pd=0.8u as=79.8f ps=0.8u w=0.42u l=0.13u
X739 a_55836_43159# VSS cap_cmim l=6.99u w=6.99u
X740 a_53774_20178# 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.sg13g2_dfrbp_1_0.CLK VDD VDD sg13_lv_pmos ad=0.34p pd=2.68u as=0.19p ps=1.38u w=1u l=0.13u
X741 VSS a_53774_20178# a_53738_20514# VSS sg13_lv_nmos ad=0.1544p pd=1.235u as=0.2516p ps=2.16u w=0.74u l=0.13u
X742 VDD a_53022_43738# a_55742_43159# VDD sg13_lv_pmos ad=59f pd=0.74u as=59.75f ps=0.745u w=0.2u l=0.13u
X743 a_45579_29803# CLK_IN a_46749_30782# VSS sg13_lv_nmos ad=79.8f pd=0.8u as=0.1428p ps=1.52u w=0.42u l=0.15u
X744 a_62119_20605# a_61887_20534# a_61394_20220# VDD sg13_lv_pmos ad=79.8f pd=0.8u as=0.1428p ps=1.52u w=0.42u l=0.13u
X745 a_62654_21971# a_61691_22290# a_62270_22299# VDD sg13_lv_pmos ad=0.17695p pd=1.56u as=0.19p ps=1.38u w=1u l=0.13u
X746 a_60479_25023# a_60385_24947# a_60385_24947# VSS sg13_lv_nmos ad=0.2307p pd=1.615u as=0.102p ps=1.28u w=0.3u l=0.13u
X747 a_64809_23027# a_64383_23628# a_64383_23300# VDD sg13_lv_pmos ad=51.45f pd=0.665u as=79.8f ps=0.8u w=0.42u l=0.13u
X748 3bit_freq_divider_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 3bit_freq_divider_0.dff_nclk_0.nCLK VSS VSS sg13_lv_nmos ad=0.259p pd=2.18u as=0.259p ps=2.18u w=0.74u l=0.13u
X749 a_64419_23654# a_64383_23628# a_64383_23889# VSS sg13_lv_nmos ad=54.6f pd=0.68u as=0.2017p ps=1.48u w=0.42u l=0.13u
X750 VSS vco_wob_0.vctl VSS VSS sg13_lv_nmos ad=0.1005p pd=1.34u as=0 ps=0 w=0.15u l=0.13u
X751 a_52886_21392# X2 VSS VSS sg13_lv_nmos ad=0.17462p pd=1.185u as=0.15245p ps=1.17u w=0.55u l=0.13u
X752 a_58536_54976# charge_pump_0.bias_n VSS VSS sg13_lv_nmos ad=0.34p pd=2.68u as=0.34p ps=2.68u w=1u l=1u
X753 VSS a_61707_25000# 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.D VSS sg13_lv_nmos ad=0.3108p pd=2.32u as=0.1628p ps=1.18u w=0.74u l=0.13u
X754 VDD a_53022_43738# a_57084_43159# VDD sg13_lv_pmos ad=59f pd=0.74u as=59.75f ps=0.745u w=0.2u l=0.13u
X755 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.nQ a_62654_21971# VDD VDD sg13_lv_pmos ad=0.7616p pd=3.6u as=0.2163p ps=1.55u w=1.12u l=0.13u
X756 VDD 3bit_freq_divider_0.sg13g2_nand2_1_0.Y 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.sg13g2_dfrbp_1_0.CLK VDD sg13_lv_pmos ad=0.392p pd=2.94u as=0.392p ps=2.94u w=1.12u l=0.13u
X757 VSS charge_pump_0.vout VSS VSS sg13_lv_nmos ad=0.285p pd=1.88u as=0 ps=0 w=1.5u l=0.65u
C0 a_52924_22885# VDD 0.20953f
C1 a_54472_22885# 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.D 0.12185f
C2 a_63463_23728# 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.Q 0.12519f
C3 3bit_freq_divider_1.dff_nclk_0.nCLK a_61394_20220# 0.37259f
C4 3bit_freq_divider_1.dff_nclk_0.nCLK a_63255_21488# 0.10313f
C5 3bit_freq_divider_1.sg13g2_or3_1_0.C 3bit_freq_divider_1.dff_nclk_0.nCLK 0.13894f
C6 a_55948_56737# charge_pump_0.bias_p 0.02673f
C7 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.Q a_61878_21130# 0.02559f
C8 3bit_freq_divider_1.sg13g2_or3_1_0.C Y1 0.16352f
C9 a_58453_40283# a_58515_40413# 0.10827f
C10 a_51684_22284# VDD 0.36995f
C11 3bit_freq_divider_0.dff_nclk_0.nCLK a_53968_20434# 0.32507f
C12 3bit_freq_divider_1.dff_nclk_0.nCLK a_64384_21091# 0.33258f
C13 VDD 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.nQ 0.18755f
C14 3bit_freq_divider_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 3bit_freq_divider_0.dff_nclk_0.D 0.17618f
C15 3bit_freq_divider_0.freq_div_cell_0.Cin 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.Q 0.22232f
C16 a_64383_23628# VDD 0.62587f
C17 3bit_freq_divider_0.dff_nclk_0.D a_51693_23426# 0.04146f
C18 a_62119_24117# a_61394_23732# 0.45825f
C19 3bit_freq_divider_0.dff_nclk_0.nCLK 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.D 0.21745f
C20 a_54427_40283# a_53022_43738# 0.18981f
C21 X0 m3_17285_2698# 0.30224f
C22 a_51693_23075# a_51648_24041# 0.03957f
C23 a_53968_20434# a_54504_20259# 0.45825f
C24 VDD a_60385_24717# 0.11381f
C25 VDD a_61691_22290# 0.68813f
C26 a_64384_21091# a_64714_21300# 0.02055f
C27 a_51684_22692# a_51685_23725# 0.04306f
C28 a_64459_24995# a_64398_24796# 0.0229f
C29 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.D a_54504_20259# 0.3562f
C30 a_63255_25000# Y0 0.39999f
C31 a_55345_24897# VDD 0.45478f
C32 VDD a_54494_43159# 1.29885f
C33 3bit_freq_divider_0.sg13g2_or3_1_0.B 3bit_freq_divider_0.sg13g2_or3_1_0.C 1.00414f
C34 a_53738_22270# a_53968_22190# 0.13068f
C35 a_53738_22270# 3bit_freq_divider_0.dff_nclk_0.nCLK 0.18642f
C36 a_51622_24863# a_51759_25014# 0.14868f
C37 a_51684_22692# X1 0.03873f
C38 a_64383_23706# VDD 0.30655f
C39 3bit_freq_divider_1.dff_nclk_0.nRST a_64384_24445# 0.04054f
C40 3bit_freq_divider_0.EN 3bit_freq_divider_1.sg13g2_nand2_1_0.Y 0.12799f
C41 a_53065_21935# a_53899_22244# 0.03957f
C42 a_57084_43159# a_57178_43159# 0.42665f
C43 X2 a_52886_21392# 0.39847f
C44 a_61887_24046# a_62119_24117# 0.13068f
C45 a_64419_23326# a_64383_23889# 0.03957f
C46 Y2 Y0 0.0326f
C47 VDD 3bit_freq_divider_0.dff_nclk_0.nRST 0.60215f
C48 3bit_freq_divider_0.freq_div_cell_0.Cout 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.Q 0.42266f
C49 m5_17331_2744# m6_17427_2840# 84.0579f
C50 a_61887_20534# a_62270_20543# 0.66077f
C51 CLK_IN m5_17331_2744# 0.42278f
C52 a_61394_21976# 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.08213f
C53 VDD a_53445_20214# 0.30479f
C54 a_64383_23628# a_64383_23706# 0.04324f
C55 a_61394_23732# VDD 0.38531f
C56 a_51684_22284# 3bit_freq_divider_0.dff_nclk_0.nRST 0.34874f
C57 VDD 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.3071f
C58 a_61691_20534# a_61394_20220# 0.17766f
C59 VDD a_63426_24642# 0.20944f
C60 a_52924_24641# a_52886_24904# 0.36535f
C61 3bit_freq_divider_1.dff_nclk_0.nCLK a_61887_20534# 0.18209f
C62 a_64383_23300# 3bit_freq_divider_1.dff_nclk_0.D 0.04146f
C63 VDD 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.D 0.9437f
C64 a_59799_40285# 3bit_freq_divider_0.CLK_IN 0.11621f
C65 VDD a_54842_49733# 0.03367f
C66 a_60967_23234# 3bit_freq_divider_1.sg13g2_nand2_1_0.Y 0.08797f
C67 a_52886_24904# 3bit_freq_divider_0.sg13g2_or3_1_0.C 0.23357f
C68 a_54472_22885# 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.Q 0.02559f
C69 a_53152_43159# a_54400_43159# 0.09188f
C70 a_64384_21091# a_64714_21414# 0.014f
C71 a_52950_22157# VDD 0.2364f
C72 3bit_freq_divider_0.dff_nclk_0.nCLK a_54504_22015# 0.37259f
C73 a_55948_56737# VDD 0.31573f
C74 a_53774_21934# 3bit_freq_divider_0.dff_nclk_0.nCLK 0.35569f
C75 a_53968_22190# a_54504_22015# 0.45825f
C76 a_53774_21934# a_53968_22190# 0.05314f
C77 a_54472_24641# 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.Q 0.02559f
C78 a_55742_43159# a_55836_43159# 0.42148f
C79 a_63463_20216# a_62654_20215# 0.09575f
C80 a_52886_21392# 3bit_freq_divider_0.sg13g2_or3_1_0.A 0.23182f
C81 X2 3bit_freq_divider_0.dff_nclk_0.nCLK 0.64366f
C82 a_60385_24947# a_60584_24580# 0.0229f
C83 CLK_IN a_48909_28913# 0.12375f
C84 a_63255_23244# 3bit_freq_divider_1.sg13g2_or3_1_0.B 0.23215f
C85 vco_wob_0.vctl a_57112_40850# 0.05026f
C86 a_56828_53480# charge_pump_0.bias_n 0.01798f
C87 VDD a_53774_20178# 0.67672f
C88 a_53445_23726# 3bit_freq_divider_0.dff_nclk_0.nCLK 0.24213f
C89 Y2 3bit_freq_divider_1.sg13g2_or3_1_0.B 0.1586f
C90 3bit_freq_divider_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK a_51631_22774# 0.33833f
C91 3bit_freq_divider_0.EN X0 0.11772f
C92 a_61887_24046# VDD 0.22153f
C93 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.Q 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.nQ 0.02712f
C94 Y1 m3_17285_2698# 0.2919f
C95 a_51631_22774# a_51693_23426# 0.05331f
C96 a_54472_22885# 3bit_freq_divider_0.freq_div_cell_0.Cin 0.01011f
C97 3bit_freq_divider_1.dff_nclk_0.nCLK a_63426_21130# 0.03449f
C98 a_62654_21971# a_63463_21972# 0.09575f
C99 a_53445_23726# a_53065_23691# 0.41048f
C100 a_53738_24026# a_53899_24000# 0.66077f
C101 a_63426_22886# a_63255_23244# 0.36535f
C102 m6_17427_2840# Y0 1.19758f
C103 3bit_freq_divider_0.dff_nclk_0.D PFD_0.VCO_CLK 0.01884f
C104 a_61675_21130# a_61707_21488# 0.0104f
C105 a_61878_24642# VDD 0.21401f
C106 VDD a_52886_21392# 0.26051f
C107 3bit_freq_divider_0.dff_nclk_0.nCLK 3bit_freq_divider_0.sg13g2_or3_1_0.A 0.48568f
C108 Y2 a_62654_21971# 0.02368f
C109 a_57178_43159# 3bit_freq_divider_0.CLK_IN 0.20831f
C110 3bit_freq_divider_1.freq_div_cell_0.Cin a_61707_25000# 0.01154f
C111 a_47954_28913# VDD 0.45155f
C112 a_52924_22885# a_52886_23148# 0.36535f
C113 VDD a_51648_24041# 0.41893f
C114 VDD a_64384_24445# 0.24105f
C115 a_52886_23148# VDD 0.25998f
C116 VDD a_52944_43077# 0.7984f
C117 a_61394_23732# 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.08213f
C118 m6_17427_2840# m7_16847_2260# 25.5177f
C119 VDD a_51600_24907# 0.04155f
C120 CLK_IN m7_16847_2260# 1.44946f
C121 a_58515_40413# a_53022_43738# 0.06975f
C122 3bit_freq_divider_0.EN 3bit_freq_divider_0.CLK_IN 0.41907f
C123 a_61691_20534# a_61887_20534# 0.45047f
C124 a_51684_22692# 3bit_freq_divider_0.sg13g2_or3_1_0.C 0.03556f
C125 3bit_freq_divider_0.freq_div_cell_1.Cout 3bit_freq_divider_0.freq_div_cell_0.Cout 0.09134f
C126 a_62270_22299# a_62654_21971# 0.03957f
C127 3bit_freq_divider_1.dff_nclk_0.nCLK a_62654_23727# 0.29516f
C128 a_52924_22885# 3bit_freq_divider_0.dff_nclk_0.nCLK 0.03415f
C129 VDD 3bit_freq_divider_1.sg13g2_nand2_1_0.Y 3.38844f
C130 m6_17427_2840# X0 1.23795f
C131 a_57311_42591# a_57178_43159# 0.22378f
C132 a_53968_22190# VDD 0.31854f
C133 3bit_freq_divider_0.dff_nclk_0.nCLK VDD 2.90191f
C134 3bit_freq_divider_1.freq_div_cell_0.Cin a_60967_24990# 0.13167f
C135 a_57173_40413# a_57112_40850# 0.03159f
C136 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.Q 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.D 0.22983f
C137 a_51622_24863# a_51721_24988# 0.0229f
C138 3bit_freq_divider_1.dff_nclk_0.nCLK a_63463_21972# 0.05956f
C139 3bit_freq_divider_1.sg13g2_tiehi_1.L_HI 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.Q 0.42892f
C140 VDD a_53058_43159# 1.37421f
C141 a_63255_25000# Y1 0.01849f
C142 Y0 VDD 0.55412f
C143 a_45451_28860# PFD_0.VCO_CLK 0.12714f
C144 a_57111_40283# a_57173_40413# 0.11922f
C145 vco_wob_0.vctl 3bit_freq_divider_0.CLK_IN 0.50349f
C146 a_53065_20179# a_53738_20514# 0.40027f
C147 a_53774_20178# a_53445_20214# 0.04324f
C148 VDD a_53065_23691# 0.44373f
C149 VDD a_57084_43159# 1.35049f
C150 a_45658_27900# PFD_0.VCO_CLK 0.17296f
C151 3bit_freq_divider_0.dff_nclk_0.nCLK 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.nQ 0.02505f
C152 3bit_freq_divider_1.dff_nclk_0.nCLK a_63255_23244# 0.10223f
C153 nEN a_56742_53480# 0.28042f
C154 a_64398_24796# CLK_OUT 0.02652f
C155 a_55831_40413# a_53022_43738# 0.04637f
C156 a_62270_24055# a_61691_24046# 0.04304f
C157 a_61887_24046# a_61394_23732# 0.47248f
C158 3bit_freq_divider_0.freq_div_cell_0.Cout 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.01369f
C159 VDD a_54504_20259# 0.36995f
C160 a_63255_25000# a_63223_24642# 0.0104f
C161 a_63255_23244# Y1 0.39563f
C162 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.D 3bit_freq_divider_0.freq_div_cell_0.Cout 0.084f
C163 Y2 3bit_freq_divider_1.dff_nclk_0.nCLK 0.86741f
C164 a_61887_24046# 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.01324f
C165 a_54434_24904# 3bit_freq_divider_0.freq_div_cell_0.Cin 0.01154f
C166 Y2 Y1 2.64011f
C167 3bit_freq_divider_1.freq_div_cell_0.Cout 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.01369f
C168 a_53065_23691# 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.nQ 0.05822f
C169 a_53774_23690# a_54504_23771# 0.17766f
C170 a_63255_21488# a_63223_21130# 0.0104f
C171 VDD a_57111_40283# 1.36202f
C172 a_53968_20434# a_53899_20488# 0.70262f
C173 a_55831_40413# a_55770_40850# 0.03778f
C174 a_55345_21385# 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.Q 0.30546f
C175 a_57311_42591# vco_wob_0.vctl 0.08436f
C176 a_51648_24041# 3bit_freq_divider_0.dff_nclk_0.nRST 0.30513f
C177 a_59800_40852# 3bit_freq_divider_0.CLK_IN 0.13041f
C178 a_55769_40283# a_55831_40413# 0.12854f
C179 3bit_freq_divider_1.dff_nclk_0.nCLK a_62270_22299# 0.17328f
C180 a_54434_23148# VDD 0.2676f
C181 3bit_freq_divider_0.dff_nclk_0.nRST a_51600_24907# 0.01267f
C182 a_62900_20179# a_62654_20215# 0.41048f
C183 a_53350_21129# a_52886_21392# 0.0104f
C184 a_56013_24979# VDD 0.11379f
C185 a_64383_23434# a_64383_23300# 0.13068f
C186 3bit_freq_divider_0.dff_nclk_0.D a_51631_22774# 0.03728f
C187 X0 VDD 1.32697f
C188 a_51622_24863# PFD_0.VCO_CLK 0.02673f
C189 a_53065_20179# 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.nQ 0.0571f
C190 a_55836_43159# a_53022_43738# 0.04103f
C191 X2 a_52924_21129# 0.02265f
C192 3bit_freq_divider_1.sg13g2_or3_1_0.B VDD 0.10974f
C193 a_62654_23727# a_63463_23728# 0.09575f
C194 3bit_freq_divider_1.freq_div_cell_0.Cin a_60967_23234# 0.13034f
C195 m5_16847_2260# m6_16847_2260# 0.13106p
C196 a_51693_23075# X1 0.01284f
C197 a_55862_56737# charge_pump_0.bias_n 0.34812f
C198 3bit_freq_divider_0.dff_nclk_0.nCLK a_53445_20214# 0.26292f
C199 a_54627_42591# vco_wob_0.vctl 0.07714f
C200 X2 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.Q 0.17317f
C201 3bit_freq_divider_1.sg13g2_nand2_1_0.Y 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.1064f
C202 3bit_freq_divider_0.EN X1 0.5347f
C203 a_63426_22886# VDD 0.20834f
C204 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.D 0.40308f
C205 3bit_freq_divider_0.sg13g2_or3_1_0.B a_51648_21103# 0.26158f
C206 a_56742_53480# charge_pump_0.bias_p 0.04781f
C207 3bit_freq_divider_0.freq_div_cell_0.Cin 3bit_freq_divider_0.sg13g2_tiehi_1.L_HI 0.14552f
C208 a_56038_24617# VDD 0.0448f
C209 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.Q a_62654_20215# 0.01984f
C210 a_62119_24117# 3bit_freq_divider_1.dff_nclk_0.nCLK 0.32742f
C211 VDD a_60967_21478# 0.45855f
C212 VDD a_62654_21971# 0.4336f
C213 3bit_freq_divider_1.sg13g2_nand2_1_0.Y 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.D 0.05067f
C214 VDD a_61707_21488# 0.2676f
C215 m6_17427_2840# Y1 1.19758f
C216 a_53147_40413# a_53022_43738# 0.08011f
C217 3bit_freq_divider_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK a_51684_22692# 0.01473f
C218 a_53152_43159# a_53022_43738# 0.08218f
C219 Y0 a_63426_24642# 0.01851f
C220 a_51684_22692# a_51693_23426# 0.13068f
C221 a_60528_49446# charge_pump_0.vout 0.01545f
C222 VDD 3bit_freq_divider_0.CLK_IN 1.60757f
C223 a_52924_21129# 3bit_freq_divider_0.sg13g2_or3_1_0.A 0.10614f
C224 3bit_freq_divider_0.freq_div_cell_1.Cout 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.D 0.04623f
C225 a_52950_22157# 3bit_freq_divider_0.dff_nclk_0.nCLK 0.05957f
C226 a_61707_23244# a_61675_22886# 0.0104f
C227 Y2 a_62900_21935# 0.0145f
C228 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.Q a_63463_20216# 0.12389f
C229 m4_17285_2698# CLK_OUT 0.3817f
C230 a_52950_20401# 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.nQ 0.21609f
C231 a_54434_24904# a_54472_24641# 0.36535f
C232 a_54489_40413# a_54428_40850# 0.03943f
C233 VDD a_55941_24882# 0.10494f
C234 a_53152_43159# a_53285_42591# 0.22378f
C235 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.nQ 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.Q 0.02712f
C236 a_53738_24026# 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.01324f
C237 vco_wob_0.vctl a_54428_40850# 0.04894f
C238 X2 X1 0.01072f
C239 3bit_freq_divider_1.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 3bit_freq_divider_1.dff_nclk_0.nCLK 0.10701f
C240 a_54427_40283# a_54489_40413# 0.12991f
C241 a_59097_54704# charge_pump_0.bias_n 0.01331f
C242 3bit_freq_divider_0.dff_nclk_0.nCLK a_53774_20178# 0.35517f
C243 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.Q 3bit_freq_divider_0.freq_div_cell_0.Cout 0.22232f
C244 a_54434_24904# 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.Q 0.46099f
C245 X0 3bit_freq_divider_0.dff_nclk_0.nRST 0.14477f
C246 a_62654_21971# a_61691_22290# 0.02302f
C247 a_62270_22299# a_61887_22290# 0.66077f
C248 3bit_freq_divider_1.freq_div_cell_0.Cout 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.Q 0.42266f
C249 a_54898_22885# a_54434_23148# 0.0104f
C250 a_52886_24904# 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.Q 0.14987f
C251 a_53968_23946# VDD 0.32286f
C252 a_64419_23326# 3bit_freq_divider_1.dff_nclk_0.D 0.01591f
C253 3bit_freq_divider_0.freq_div_cell_0.Cout a_54434_21392# 0.12082f
C254 VDD a_62270_20543# 0.24492f
C255 3bit_freq_divider_1.dff_nclk_0.nCLK 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.nQ 0.08552f
C256 m5_17331_2744# Y0 0.40842f
C257 VDD a_52924_21129# 0.20953f
C258 a_55345_21385# 3bit_freq_divider_0.freq_div_cell_1.Cout 0.13166f
C259 a_53774_20178# a_54504_20259# 0.17766f
C260 3bit_freq_divider_0.EN 3bit_freq_divider_0.freq_div_cell_1.Cout 0.01552f
C261 a_51648_24438# VDD 0.24104f
C262 a_47954_28913# a_48909_28913# 0.39061f
C263 a_46817_27899# PFD_0.VCO_CLK 0.92547f
C264 3bit_freq_divider_1.sg13g2_or3_1_0.C a_64419_23326# 0.01089f
C265 3bit_freq_divider_0.dff_nclk_0.nCLK a_52886_21392# 0.10313f
C266 3bit_freq_divider_1.dff_nclk_0.nCLK VDD 2.89514f
C267 a_64383_23300# 3bit_freq_divider_1.dff_nclk_0.nRST 0.31482f
C268 VDD Y1 0.44908f
C269 charge_pump_0.bias_p charge_pump_0.vout 0.02402f
C270 nEN charge_pump_0.bias_n 0.06869f
C271 VDD a_60584_24580# 0.10495f
C272 3bit_freq_divider_0.freq_div_cell_0.Cout 3bit_freq_divider_0.freq_div_cell_0.Cin 0.10559f
C273 VDD 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.Q 1.42261f
C274 3bit_freq_divider_1.freq_div_cell_0.Cin VDD 1.21632f
C275 a_52886_23148# 3bit_freq_divider_0.dff_nclk_0.nCLK 0.10223f
C276 vco_wob_0.vctl charge_pump_0.vout 0.05724f
C277 a_59799_40285# a_58515_40413# 0.46077f
C278 a_52950_23913# 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.Q 0.12519f
C279 a_53738_22270# 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.01324f
C280 a_54627_42591# VDD 0.01623f
C281 a_52944_43077# a_53058_43159# 0.08875f
C282 a_62270_22299# a_62119_22361# 0.70262f
C283 PFD_0.DOWN CLK_IN 0.06328f
C284 a_54472_24641# 3bit_freq_divider_0.sg13g2_tiehi_1.L_HI 0.01011f
C285 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.nQ VDD 0.18275f
C286 PFD_0.DOWN a_54357_49278# 0.04759f
C287 VDD a_64714_21300# 0.01263f
C288 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.D VDD 0.97883f
C289 3bit_freq_divider_1.dff_nclk_0.nCLK a_61691_22290# 0.35569f
C290 m5_17331_2744# X0 0.42278f
C291 3bit_freq_divider_0.freq_div_cell_0.Cout 3bit_freq_divider_0.sg13g2_nand2_1_0.Y 0.3426f
C292 a_51693_23075# 3bit_freq_divider_0.sg13g2_or3_1_0.C 0.01089f
C293 a_51685_23725# VDD 0.30547f
C294 a_61707_21488# 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.D 0.24715f
C295 a_45658_27900# a_46817_27899# 0.43194f
C296 a_55969_42591# a_55836_43159# 0.22378f
C297 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.Q 3bit_freq_divider_0.sg13g2_tiehi_1.L_HI 0.42892f
C298 a_62900_23691# 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.nQ 0.10118f
C299 a_53968_22190# 3bit_freq_divider_0.dff_nclk_0.nCLK 0.32534f
C300 a_60385_24717# a_60584_24580# 0.14868f
C301 3bit_freq_divider_0.freq_div_cell_0.Cout a_54472_21129# 0.01011f
C302 a_64424_22200# 3bit_freq_divider_1.dff_nclk_0.D 0.43097f
C303 a_52924_22885# X1 0.02265f
C304 3bit_freq_divider_1.dff_nclk_0.D a_64383_23889# 0.09445f
C305 a_53022_43738# a_54400_43159# 0.19723f
C306 VDD X1 1.47452f
C307 a_54357_49278# charge_pump_0.vout 0.01432f
C308 3bit_freq_divider_0.dff_nclk_0.nCLK a_53065_23691# 0.29533f
C309 3bit_freq_divider_0.EN charge_pump_0.bias_n 0.02661f
C310 VDD a_53899_20488# 0.24492f
C311 3bit_freq_divider_0.dff_nclk_0.nCLK a_54504_20259# 0.37259f
C312 VDD a_54428_40850# 0.01457f
C313 a_54504_22015# 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.08213f
C314 a_51684_22284# X1 0.0269f
C315 a_53774_21934# 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.33731f
C316 a_51684_22692# 3bit_freq_divider_0.dff_nclk_0.D 0.0175f
C317 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.D a_54504_22015# 0.3562f
C318 X0 a_51648_24041# 0.0271f
C319 a_53774_21934# 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.D 0.01446f
C320 a_51648_24438# 3bit_freq_divider_0.dff_nclk_0.nRST 0.04054f
C321 a_53774_23690# a_53899_24000# 0.04304f
C322 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.D a_61691_22290# 0.01446f
C323 a_46749_30782# a_47777_29803# 0.4544f
C324 VDD a_54427_40283# 1.36925f
C325 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.Q a_62654_23727# 0.0119f
C326 charge_pump_0.bias_n charge_pump_0.bias_p 1.09436f
C327 a_63463_23728# VDD 0.2349f
C328 a_54627_42591# a_54494_43159# 0.22378f
C329 a_58453_40283# a_53022_43738# 0.19288f
C330 a_61707_25000# 3bit_freq_divider_1.sg13g2_tiehi_1.L_HI 0.12082f
C331 PFD_0.DOWN VDD 1.56226f
C332 3bit_freq_divider_1.dff_nclk_0.nCLK a_61394_23732# 0.37259f
C333 VDD a_61887_22290# 0.21577f
C334 VDD a_61691_20534# 0.67211f
C335 3bit_freq_divider_1.dff_nclk_0.nCLK 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.60301f
C336 Y0 m7_16847_2260# 1.40976f
C337 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.Q a_63463_21972# 0.12389f
C338 3bit_freq_divider_0.freq_div_cell_0.Cin 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.01369f
C339 X2 3bit_freq_divider_0.sg13g2_or3_1_0.C 0.04643f
C340 VDD a_62900_21935# 0.30801f
C341 3bit_freq_divider_0.freq_div_cell_0.Cin 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.D 0.084f
C342 a_63426_24642# Y1 0.01474f
C343 a_53350_22885# a_52886_23148# 0.0104f
C344 3bit_freq_divider_1.dff_nclk_0.nCLK 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.D 0.21745f
C345 3bit_freq_divider_1.freq_div_cell_0.Cin 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.01369f
C346 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.sg13g2_dfrbp_1_0.CLK VDD 0.27798f
C347 a_55742_43159# a_53022_43738# 0.19603f
C348 a_63255_23244# 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.Q 0.12248f
C349 VDD a_61878_21130# 0.21321f
C350 CLK_IN a_47777_29803# 0.17902f
C351 a_54434_21392# 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.D 0.24715f
C352 a_64383_23300# VDD 0.29403f
C353 VDD charge_pump_0.vout 0.06128f
C354 Y2 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.Q 0.20327f
C355 3bit_freq_divider_0.EN a_58536_54976# 0.21462f
C356 a_53445_23726# a_53738_24026# 0.04306f
C357 a_45579_29803# a_46749_30782# 0.25388f
C358 3bit_freq_divider_1.sg13g2_tiehi_1.L_HI a_60967_24990# 0.21784f
C359 a_51685_23725# 3bit_freq_divider_0.dff_nclk_0.nRST 0.25925f
C360 a_53147_40413# a_53085_40283# 0.10818f
C361 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 3bit_freq_divider_0.sg13g2_nand2_1_0.Y 0.1064f
C362 3bit_freq_divider_0.freq_div_cell_1.Cout VDD 0.4595f
C363 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.D 3bit_freq_divider_0.sg13g2_nand2_1_0.Y 0.04726f
C364 a_58515_40413# vco_wob_0.vctl 0.02267f
C365 a_61691_22290# a_61887_22290# 0.45047f
C366 a_64383_23628# a_64383_23300# 0.05314f
C367 a_61887_20534# a_62654_20215# 0.40027f
C368 a_61878_22886# VDD 0.21321f
C369 3bit_freq_divider_1.freq_div_cell_0.Cout 3bit_freq_divider_1.freq_div_cell_1.Cout 0.09134f
C370 a_58454_40850# vco_wob_0.vctl 0.04998f
C371 3bit_freq_divider_0.dff_nclk_0.nRST X1 0.08188f
C372 a_61691_24046# 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.D 0.01446f
C373 a_58536_54976# charge_pump_0.bias_p 0.38944f
C374 a_61691_22290# a_62900_21935# 0.04324f
C375 a_60967_21478# 3bit_freq_divider_1.sg13g2_nand2_1_0.Y 0.08797f
C376 a_61887_24046# 3bit_freq_divider_1.dff_nclk_0.nCLK 0.18489f
C377 X0 m7_16847_2260# 1.44946f
C378 VDD a_62119_22361# 0.31854f
C379 a_52950_22157# 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.nQ 0.21609f
C380 a_64383_23434# a_64419_23326# 0.66077f
C381 m5_17331_2744# Y1 0.40842f
C382 a_63255_21488# 3bit_freq_divider_1.sg13g2_or3_1_0.A 0.23182f
C383 a_53738_20514# a_53968_20434# 0.13068f
C384 CLK_IN a_45579_29803# 1.21724f
C385 3bit_freq_divider_1.sg13g2_nand2_1_0.Y 3bit_freq_divider_0.CLK_IN 0.2618f
C386 a_51708_21299# a_51648_21103# 0.02055f
C387 a_60967_23234# 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.Q 0.30546f
C388 a_52924_21129# a_52886_21392# 0.36535f
C389 3bit_freq_divider_1.sg13g2_or3_1_0.A a_64384_21091# 0.31317f
C390 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK VDD 0.29872f
C391 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.D VDD 0.97883f
C392 a_54489_40413# a_55831_40413# 0.72984f
C393 a_59800_40852# a_58515_40413# 0.21632f
C394 VDD a_47777_29803# 1.07957f
C395 a_52950_20401# a_53065_20179# 0.09575f
C396 a_51693_23075# a_51693_23426# 0.70262f
C397 a_53147_40413# a_53086_40850# 0.04971f
C398 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.D 3bit_freq_divider_0.sg13g2_nand2_1_0.Y 0.05067f
C399 VDD a_52924_24641# 0.21522f
C400 a_51648_24438# a_51648_24041# 0.09575f
C401 a_55836_43159# a_57178_43159# 0.91818f
C402 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.Q a_52886_21392# 0.12248f
C403 a_55831_40413# vco_wob_0.vctl 0.04109f
C404 a_62900_23691# a_61691_24046# 0.04324f
C405 a_53445_21970# a_53738_22270# 0.04306f
C406 a_54434_21392# a_54898_21129# 0.0104f
C407 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.D a_54472_21129# 0.12185f
C408 VDD 3bit_freq_divider_0.sg13g2_or3_1_0.C 0.20391f
C409 3bit_freq_divider_0.EN a_58734_56203# 0.07729f
C410 a_62119_22361# a_61691_22290# 0.05314f
C411 a_53738_24026# VDD 0.22151f
C412 a_53968_23946# 3bit_freq_divider_0.dff_nclk_0.nCLK 0.32517f
C413 VDD charge_pump_0.bias_n 0.83592f
C414 a_51684_22692# a_51631_22774# 0.45006f
C415 a_56038_24617# a_56013_24979# 0.01952f
C416 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.D a_61691_20534# 0.01446f
C417 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.D a_54472_24641# 0.12185f
C418 3bit_freq_divider_0.dff_nclk_0.nCLK a_52924_21129# 0.03449f
C419 a_53774_20178# a_53899_20488# 0.04304f
C420 charge_pump_0.bias_p a_58734_56203# 0.03822f
C421 a_63426_22886# 3bit_freq_divider_1.sg13g2_or3_1_0.B 0.10697f
C422 a_57173_40413# a_58515_40413# 0.58365f
C423 3bit_freq_divider_1.dff_nclk_0.nCLK 3bit_freq_divider_1.sg13g2_nand2_1_0.Y 0.23907f
C424 a_58454_40850# a_57173_40413# 0.22936f
C425 VDD a_45579_29803# 0.45874f
C426 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.D 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.Q 0.22983f
C427 a_61878_21130# 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.D 0.12185f
C428 3bit_freq_divider_1.dff_nclk_0.D CLK_OUT 0.01884f
C429 a_64383_23434# a_64424_22200# 0.47248f
C430 a_55345_21385# 3bit_freq_divider_0.sg13g2_nand2_1_0.Y 0.08797f
C431 VDD a_56137_24678# 0.11858f
C432 a_64383_23434# a_64383_23889# 0.40027f
C433 3bit_freq_divider_1.freq_div_cell_0.Cin 3bit_freq_divider_1.sg13g2_nand2_1_0.Y 0.25573f
C434 3bit_freq_divider_0.EN 3bit_freq_divider_0.sg13g2_nand2_1_0.Y 0.12847f
C435 a_51685_23725# a_51648_24041# 0.41048f
C436 3bit_freq_divider_0.dff_nclk_0.nCLK 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.Q 1.0402f
C437 a_55836_43159# vco_wob_0.vctl 0.02497f
C438 charge_pump_0.vout a_54842_49733# 0.02265f
C439 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.D 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.Q 0.22983f
C440 Y0 Y1 1.97044f
C441 a_62270_24055# a_62654_23727# 0.03957f
C442 a_53065_21935# a_53738_22270# 0.40027f
C443 a_53774_21934# a_53445_21970# 0.04324f
C444 a_56013_24979# a_55941_24882# 0.14868f
C445 m4_17285_2698# m3_17285_2698# 0.20496p
C446 a_58426_43159# a_53022_43738# 0.10045f
C447 VDD a_58515_40413# 1.36426f
C448 a_52886_23148# X1 0.39847f
C449 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.nQ 3bit_freq_divider_0.dff_nclk_0.nCLK 0.08742f
C450 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.sg13g2_dfrbp_1_0.CLK a_53774_20178# 0.33731f
C451 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.D 3bit_freq_divider_1.sg13g2_nand2_1_0.Y 0.05125f
C452 a_61707_23244# VDD 0.2676f
C453 a_61394_20220# a_62119_20605# 0.45825f
C454 VDD a_51759_25014# 0.0834f
C455 VDD a_58536_54976# 0.98046f
C456 a_64398_24796# 3bit_freq_divider_1.dff_nclk_0.nRST 0.10221f
C457 a_55831_40413# a_57173_40413# 0.7336f
C458 a_55345_23141# 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.Q 0.30546f
C459 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.sg13g2_dfrbp_1_0.CLK a_61394_20220# 0.08213f
C460 a_62654_23727# 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.nQ 0.05822f
C461 m7_16847_2260# Y1 1.40976f
C462 a_53147_40413# a_54489_40413# 0.35714f
C463 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.Q a_63255_21488# 0.12248f
C464 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.Q VDD 1.41895f
C465 a_64419_23326# 3bit_freq_divider_1.dff_nclk_0.nRST 0.16457f
C466 a_53774_23690# 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.33731f
C467 a_53147_40413# vco_wob_0.vctl 0.04038f
C468 a_53152_43159# vco_wob_0.vctl 0.02282f
C469 3bit_freq_divider_0.dff_nclk_0.nRST 3bit_freq_divider_0.sg13g2_or3_1_0.C 0.57774f
C470 a_54504_23771# 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.08213f
C471 a_54434_24904# 3bit_freq_divider_0.sg13g2_tiehi_1.L_HI 0.12082f
C472 3bit_freq_divider_0.dff_nclk_0.nCLK X1 0.26228f
C473 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.D a_53774_23690# 0.01446f
C474 a_51648_24438# X0 0.01187f
C475 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.D a_54504_23771# 0.3562f
C476 3bit_freq_divider_1.sg13g2_or3_1_0.C 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.Q 0.05745f
C477 VDD a_55831_40413# 1.08631f
C478 3bit_freq_divider_0.dff_nclk_0.nCLK a_53899_20488# 0.17248f
C479 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.Q a_52924_22885# 0.01011f
C480 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.Q VDD 1.42273f
C481 3bit_freq_divider_1.dff_nclk_0.nCLK 3bit_freq_divider_1.sg13g2_or3_1_0.B 0.58488f
C482 a_53738_22270# a_53899_22244# 0.66077f
C483 a_53065_21935# a_53774_21934# 0.02335f
C484 3bit_freq_divider_1.sg13g2_or3_1_0.B Y1 0.13266f
C485 a_53285_42591# a_53022_43738# 0.02036f
C486 Y2 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.nQ 0.04535f
C487 a_55345_23141# 3bit_freq_divider_0.freq_div_cell_0.Cin 0.13034f
C488 VDD a_54434_21392# 0.2676f
C489 a_55769_40283# a_53022_43738# 0.19098f
C490 3bit_freq_divider_1.sg13g2_or3_1_0.A a_63426_21130# 0.10614f
C491 a_51693_23075# 3bit_freq_divider_0.dff_nclk_0.D 0.01591f
C492 VDD 3bit_freq_divider_1.sg13g2_tiehi_1.L_HI 0.7718f
C493 VDD a_61394_21976# 0.38024f
C494 3bit_freq_divider_1.dff_nclk_0.nCLK a_63426_22886# 0.03415f
C495 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.Q 3bit_freq_divider_1.freq_div_cell_1.Cout 0.2223f
C496 a_62900_20179# a_61887_20534# 0.04306f
C497 a_63426_22886# Y1 0.01971f
C498 3bit_freq_divider_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK VDD 0.28742f
C499 VDD a_51693_23426# 0.29403f
C500 3bit_freq_divider_1.dff_nclk_0.nCLK a_62654_21971# 0.31887f
C501 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 3bit_freq_divider_0.dff_nclk_0.nCLK 0.60301f
C502 VDD a_58734_56203# 0.35557f
C503 a_51685_23725# X0 0.02143f
C504 3bit_freq_divider_0.freq_div_cell_0.Cin VDD 1.21627f
C505 a_55345_23141# 3bit_freq_divider_0.sg13g2_nand2_1_0.Y 0.08797f
C506 a_51684_22284# 3bit_freq_divider_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.0838f
C507 VDD a_55836_43159# 1.00781f
C508 a_53445_21970# VDD 0.30838f
C509 a_51684_22284# a_51693_23426# 0.45825f
C510 3bit_freq_divider_0.dff_nclk_0.nRST a_51759_25014# 0.03098f
C511 a_64424_22200# 3bit_freq_divider_1.dff_nclk_0.nRST 0.34882f
C512 3bit_freq_divider_1.dff_nclk_0.nRST a_64383_23889# 0.30513f
C513 a_64398_24796# a_64362_24865# 0.14868f
C514 X0 X1 0.55463f
C515 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.Q 3bit_freq_divider_0.CLK_IN 0.02001f
C516 a_53774_21934# a_53899_22244# 0.04304f
C517 a_62270_24055# a_62119_24117# 0.70262f
C518 a_60385_24717# 3bit_freq_divider_1.sg13g2_tiehi_1.L_HI 0.02161f
C519 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.sg13g2_dfrbp_1_0.CLK a_54504_20259# 0.08213f
C520 a_61691_22290# a_61394_21976# 0.17766f
C521 a_61887_20534# a_62119_20605# 0.13068f
C522 VDD a_53738_20514# 0.19386f
C523 VDD 3bit_freq_divider_0.sg13g2_nand2_1_0.Y 3.38843f
C524 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.sg13g2_dfrbp_1_0.CLK a_61887_20534# 0.01324f
C525 VDD a_54472_21129# 0.21321f
C526 a_60967_23234# 3bit_freq_divider_1.freq_div_cell_0.Cout 0.13167f
C527 CLK_IN PFD_0.UP 0.15472f
C528 VDD a_64398_24796# 0.09559f
C529 3bit_freq_divider_1.dff_nclk_0.nCLK a_62270_20543# 0.17248f
C530 a_54357_49278# PFD_0.UP 0.30851f
C531 VDD a_53147_40413# 0.81739f
C532 CLK_OUT m3_17285_2698# 0.2919f
C533 VDD a_53152_43159# 1.05457f
C534 a_64419_23326# VDD 0.2446f
C535 3bit_freq_divider_1.sg13g2_or3_1_0.C a_64384_21091# 0.25034f
C536 a_55345_24897# 3bit_freq_divider_0.freq_div_cell_0.Cin 0.13167f
C537 3bit_freq_divider_0.dff_nclk_0.nCLK 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.60301f
C538 a_53065_21935# VDD 0.43552f
C539 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.D 3bit_freq_divider_0.dff_nclk_0.nCLK 0.21745f
C540 a_52924_21129# 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.Q 0.01011f
C541 a_51648_21103# 3bit_freq_divider_0.sg13g2_or3_1_0.A 0.31317f
C542 3bit_freq_divider_1.dff_nclk_0.nCLK Y1 0.23798f
C543 a_54494_43159# a_55836_43159# 0.88103f
C544 Y2 3bit_freq_divider_1.sg13g2_or3_1_0.A 0.10441f
C545 a_62654_23727# a_61691_24046# 0.02302f
C546 3bit_freq_divider_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 3bit_freq_divider_0.dff_nclk_0.nRST 0.16209f
C547 3bit_freq_divider_1.freq_div_cell_0.Cin 3bit_freq_divider_1.dff_nclk_0.nCLK 0.32366f
C548 a_64419_23326# a_64383_23628# 0.04304f
C549 VDD a_51721_24988# 0.08543f
C550 3bit_freq_divider_0.dff_nclk_0.nCLK 3bit_freq_divider_0.sg13g2_or3_1_0.C 0.13894f
C551 3bit_freq_divider_0.dff_nclk_0.nRST a_51693_23426# 0.3148f
C552 a_64459_24995# a_64362_24865# 0.10864f
C553 a_52950_22157# 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.Q 0.12389f
C554 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.nQ a_62654_20215# 0.0571f
C555 VDD 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.nQ 0.18065f
C556 a_53738_24026# 3bit_freq_divider_0.dff_nclk_0.nCLK 0.18638f
C557 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.Q a_63426_21130# 0.01011f
C558 a_62270_24055# VDD 0.26494f
C559 a_62654_21971# a_61887_22290# 0.40027f
C560 CLK_IN m4_17285_2698# 0.39515f
C561 a_64424_22200# 3bit_freq_divider_1.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.0838f
C562 VDD a_62654_20215# 0.42601f
C563 a_62654_21971# a_62900_21935# 0.41048f
C564 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.D 3bit_freq_divider_1.dff_nclk_0.nCLK 0.21745f
C565 a_53445_23726# a_53774_23690# 0.04324f
C566 a_53738_24026# a_53065_23691# 0.40027f
C567 VDD a_54472_24641# 0.214f
C568 VDD PFD_0.UP 0.82664f
C569 a_61675_24642# a_61707_25000# 0.0104f
C570 a_51693_23075# a_51631_22774# 0.04255f
C571 a_61878_21130# a_61707_21488# 0.36535f
C572 a_64459_24995# VDD 0.08543f
C573 VDD a_51648_21103# 0.34051f
C574 a_53152_43159# a_54494_43159# 0.77984f
C575 a_63463_20216# 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.nQ 0.21609f
C576 VDD 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.nQ 0.18204f
C577 a_53899_22244# VDD 0.26052f
C578 VDD 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.Q 1.68952f
C579 a_53445_20214# a_53738_20514# 0.04306f
C580 a_61707_25000# 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.Q 0.46099f
C581 a_51600_24907# a_51759_25014# 0.01952f
C582 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.D a_54434_23148# 0.24715f
C583 a_54434_24904# 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.D 0.24715f
C584 CLK_IN a_45451_28860# 0.13923f
C585 VDD 3bit_freq_divider_0.dff_nclk_0.D 0.84532f
C586 a_64424_22200# VDD 0.36995f
C587 VDD a_63463_20216# 0.2331f
C588 VDD a_64383_23889# 0.41974f
C589 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.nQ 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.Q 0.02712f
C590 X0 a_52924_24641# 0.02265f
C591 a_53085_40283# a_53022_43738# 0.23019f
C592 a_51684_22284# 3bit_freq_divider_0.dff_nclk_0.D 0.43097f
C593 VDD PFD_0.VCO_CLK 1.82327f
C594 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.nQ a_63463_21972# 0.21609f
C595 a_61691_20534# a_62270_20543# 0.04304f
C596 a_61394_20220# a_61887_20534# 0.47248f
C597 CLK_IN m1_17285_2698# 0.01061f
C598 3bit_freq_divider_1.freq_div_cell_0.Cout VDD 1.22849f
C599 X0 3bit_freq_divider_0.sg13g2_or3_1_0.C 0.41386f
C600 a_64424_22200# a_64383_23628# 0.17766f
C601 a_64383_23628# a_64383_23889# 0.02302f
C602 a_61878_24642# 3bit_freq_divider_1.sg13g2_tiehi_1.L_HI 0.01011f
C603 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.Q a_52886_23148# 0.12248f
C604 a_60967_24990# 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.Q 0.30546f
C605 a_63463_23728# Y1 0.03561f
C606 a_59799_40285# a_53022_43738# 0.19389f
C607 a_58653_42591# a_57178_43159# 0.03205f
C608 3bit_freq_divider_1.dff_nclk_0.nCLK a_61887_22290# 0.18493f
C609 a_62654_23727# 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.Q 0.02071f
C610 3bit_freq_divider_1.dff_nclk_0.nCLK a_61691_20534# 0.35517f
C611 a_61707_25000# 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.D 0.24715f
C612 Y2 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.nQ 0.04365f
C613 3bit_freq_divider_1.dff_nclk_0.nCLK a_62900_21935# 0.27425f
C614 VDD a_54400_43159# 1.37065f
C615 a_63255_25000# 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.Q 0.14987f
C616 a_58453_40283# a_57173_40413# 0.46167f
C617 a_56013_24979# a_56137_24678# 0.10864f
C618 a_53774_20178# a_53738_20514# 0.44698f
C619 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.nQ a_53445_20214# 0.10118f
C620 VDD a_53774_23690# 0.70098f
C621 VDD a_54504_23771# 0.38531f
C622 m2_17285_2698# m1_17285_2698# 0.20496p
C623 a_55345_24897# 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.Q 0.30546f
C624 Y2 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.Q 0.15836f
C625 3bit_freq_divider_1.dff_nclk_0.nRST CLK_OUT 0.07748f
C626 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.Q 3bit_freq_divider_0.dff_nclk_0.nCLK 1.03924f
C627 nEN a_56828_53480# 0.06208f
C628 a_52950_22157# a_53065_21935# 0.09575f
C629 a_53086_40850# a_53022_43738# 0.06371f
C630 a_62119_24117# a_61691_24046# 0.05314f
C631 VDD a_45451_28860# 0.05543f
C632 a_64383_23434# 3bit_freq_divider_1.dff_nclk_0.D 0.0175f
C633 a_45658_27900# VDD 1.00659f
C634 Y2 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.Q 0.21293f
C635 a_63255_21488# a_63426_21130# 0.36535f
C636 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.Q a_53065_23691# 0.0119f
C637 a_58426_43159# a_57178_43159# 0.1057f
C638 VDD a_58453_40283# 1.38336f
C639 a_64383_23706# a_64383_23889# 0.41048f
C640 a_64383_23434# 3bit_freq_divider_1.sg13g2_or3_1_0.C 0.03556f
C641 3bit_freq_divider_0.freq_div_cell_1.Cout 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.Q 0.2223f
C642 a_55831_40413# a_57112_40850# 0.23035f
C643 VDD 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.29872f
C644 PFD_0.DOWN a_54747_49259# 0.01456f
C645 a_58653_42591# vco_wob_0.vctl 0.08336f
C646 3bit_freq_divider_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 3bit_freq_divider_0.dff_nclk_0.nCLK 0.10701f
C647 3bit_freq_divider_0.dff_nclk_0.D 3bit_freq_divider_0.dff_nclk_0.nRST 0.76289f
C648 X2 3bit_freq_divider_0.sg13g2_or3_1_0.B 0.33008f
C649 a_57111_40283# a_55831_40413# 0.45955f
C650 3bit_freq_divider_1.dff_nclk_0.nCLK a_62119_22361# 0.32758f
C651 VDD 3bit_freq_divider_1.sg13g2_or3_1_0.A 0.12797f
C652 3bit_freq_divider_1.freq_div_cell_0.Cin a_61878_22886# 0.01011f
C653 3bit_freq_divider_0.dff_nclk_0.nCLK 3bit_freq_divider_0.freq_div_cell_0.Cin 0.32366f
C654 a_56039_25022# VDD 0.01215f
C655 VDD a_55742_43159# 1.36686f
C656 a_53445_21970# 3bit_freq_divider_0.dff_nclk_0.nCLK 0.27428f
C657 3bit_freq_divider_0.dff_nclk_0.nRST PFD_0.VCO_CLK 0.06912f
C658 m6_17427_2840# CLK_OUT 1.19758f
C659 a_54494_43159# a_54400_43159# 0.42202f
C660 a_57178_43159# a_53022_43738# 0.04298f
C661 charge_pump_0.vout a_54747_49259# 0.13589f
C662 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.Q a_54434_23148# 0.46099f
C663 a_53147_40413# a_52944_43077# 0.40206f
C664 a_62654_23727# a_62900_23691# 0.41048f
C665 a_61887_24046# a_62270_24055# 0.66077f
C666 a_53738_24026# a_53968_23946# 0.13068f
C667 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.D a_61878_22886# 0.12185f
C668 a_57084_43159# a_55836_43159# 0.09926f
C669 a_52944_43077# a_53152_43159# 0.3548f
C670 VDD a_51622_24863# 0.09559f
C671 a_58515_40413# 3bit_freq_divider_0.CLK_IN 0.83094f
C672 a_61691_22290# 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.33731f
C673 3bit_freq_divider_0.dff_nclk_0.nCLK a_53738_20514# 0.18358f
C674 a_55941_24882# a_56137_24678# 0.0229f
C675 3bit_freq_divider_0.dff_nclk_0.nCLK 3bit_freq_divider_0.sg13g2_nand2_1_0.Y 0.23907f
C676 a_54472_22885# VDD 0.21321f
C677 a_63426_22886# 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.Q 0.01011f
C678 a_61691_24046# VDD 0.69635f
C679 a_58454_40850# 3bit_freq_divider_0.CLK_IN 0.02056f
C680 VDD a_51631_22774# 0.62631f
C681 3bit_freq_divider_0.sg13g2_or3_1_0.B 3bit_freq_divider_0.sg13g2_or3_1_0.A 0.72102f
C682 a_63255_25000# 3bit_freq_divider_1.sg13g2_or3_1_0.C 0.23357f
C683 a_61887_22290# a_62900_21935# 0.04306f
C684 m6_60810_42209# a_57178_43159# 0.08511f
C685 a_60385_24558# VDD 0.04481f
C686 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.Q a_62654_21971# 0.01984f
C687 a_62900_20179# 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.nQ 0.10118f
C688 a_51684_22284# a_51631_22774# 0.17766f
C689 a_54489_40413# a_53022_43738# 0.05403f
C690 a_53152_43159# a_53058_43159# 0.42803f
C691 a_53738_20514# a_54504_20259# 0.47248f
C692 Y2 a_62900_23691# 0.01917f
C693 a_54434_23148# 3bit_freq_divider_0.freq_div_cell_0.Cin 0.12082f
C694 vco_wob_0.vctl a_53022_43738# 0.09057f
C695 a_53065_21935# 3bit_freq_divider_0.dff_nclk_0.nCLK 0.31904f
C696 VDD a_62900_20179# 0.30479f
C697 a_55742_43159# a_54494_43159# 0.10275f
C698 Y2 a_63255_21488# 0.39947f
C699 a_51684_22692# a_51693_23075# 0.66077f
C700 a_54434_24904# a_54898_24641# 0.0104f
C701 VDD CLK_OUT 0.38178f
C702 a_54489_40413# a_55770_40850# 0.23444f
C703 VDD a_60479_25023# 0.01215f
C704 a_52924_22885# 3bit_freq_divider_0.sg13g2_or3_1_0.B 0.10697f
C705 a_56742_53480# charge_pump_0.bias_n 0.05592f
C706 vco_wob_0.vctl a_55770_40850# 0.05041f
C707 VDD a_53065_20179# 0.42601f
C708 3bit_freq_divider_0.dff_nclk_0.nCLK 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.nQ 0.08555f
C709 3bit_freq_divider_0.sg13g2_or3_1_0.B VDD 0.11082f
C710 vco_wob_0.vctl a_53285_42591# 0.08086f
C711 a_60385_24558# a_60385_24717# 0.01952f
C712 a_55769_40283# a_54489_40413# 0.45379f
C713 3bit_freq_divider_1.dff_nclk_0.nRST 3bit_freq_divider_1.dff_nclk_0.D 0.7629f
C714 m4_17285_2698# m5_17331_2744# 0.1814p
C715 a_62119_22361# a_61887_22290# 0.13068f
C716 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.Q 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.nQ 0.02712f
C717 VDD 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.nQ 0.18067f
C718 a_51648_24041# 3bit_freq_divider_0.dff_nclk_0.D 0.09445f
C719 3bit_freq_divider_0.sg13g2_or3_1_0.C X1 0.20623f
C720 m6_60810_42209# vco_wob_0.vctl 0.05504f
C721 VDD a_62119_20605# 0.2982f
C722 a_59800_40852# a_53022_43738# 0.01439f
C723 a_64384_24445# a_64383_23889# 0.09575f
C724 3bit_freq_divider_1.sg13g2_or3_1_0.C 3bit_freq_divider_1.dff_nclk_0.nRST 0.57774f
C725 VDD 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.27798f
C726 a_63223_22886# a_63255_23244# 0.0104f
C727 VDD 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.Q 1.4225f
C728 a_51622_24863# 3bit_freq_divider_0.dff_nclk_0.nRST 0.10221f
C729 a_47954_28913# PFD_0.VCO_CLK 1.24436f
C730 m3_16847_2260# m4_16847_2260# 0.2063p
C731 3bit_freq_divider_1.dff_nclk_0.nCLK 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.Q 1.03922f
C732 3bit_freq_divider_1.freq_div_cell_0.Cin a_61707_23244# 0.12082f
C733 3bit_freq_divider_0.dff_nclk_0.nCLK a_51648_21103# 0.33244f
C734 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.Q Y1 0.15164f
C735 a_53899_22244# 3bit_freq_divider_0.dff_nclk_0.nCLK 0.17328f
C736 a_53968_22190# a_53899_22244# 0.70262f
C737 3bit_freq_divider_0.dff_nclk_0.nCLK 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.Q 0.08441f
C738 3bit_freq_divider_0.dff_nclk_0.nRST a_51631_22774# 0.3267f
C739 VDD 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.Q 1.66358f
C740 3bit_freq_divider_1.freq_div_cell_0.Cin 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.Q 0.42266f
C741 a_46817_27899# VDD 1.02029f
C742 a_48909_28913# PFD_0.VCO_CLK 0.1514f
C743 3bit_freq_divider_0.dff_nclk_0.nCLK 3bit_freq_divider_0.dff_nclk_0.D 0.04354f
C744 a_54434_24904# VDD 0.27564f
C745 a_61691_24046# a_61394_23732# 0.17766f
C746 VDD a_58426_43159# 1.36969f
C747 3bit_freq_divider_0.EN 3bit_freq_divider_1.freq_div_cell_1.Cout 0.01552f
C748 a_61691_24046# 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.33731f
C749 m6_16847_2260# m7_16847_2260# 39.787f
C750 VDD a_52886_24904# 0.28115f
C751 a_53065_23691# 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.Q 0.02071f
C752 PFD_0.DOWN charge_pump_0.bias_n 0.01578f
C753 a_61707_23244# 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.D 0.24715f
C754 a_57173_40413# a_53022_43738# 0.04406f
C755 a_55345_21385# 3bit_freq_divider_0.freq_div_cell_0.Cout 0.13034f
C756 3bit_freq_divider_1.freq_div_cell_0.Cout 3bit_freq_divider_1.sg13g2_nand2_1_0.Y 0.3426f
C757 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.D 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.40308f
C758 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.D 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.Q 0.22983f
C759 VDD a_52950_20401# 0.2331f
C760 3bit_freq_divider_0.sg13g2_nand2_1_0.Y 3bit_freq_divider_0.CLK_IN 0.2618f
C761 3bit_freq_divider_1.dff_nclk_0.nCLK a_61394_21976# 0.37259f
C762 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.Q a_54434_21392# 0.46099f
C763 a_57311_42591# a_55836_43159# 0.03153f
C764 charge_pump_0.bias_n charge_pump_0.vout 0.23558f
C765 VDD 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.D 0.97083f
C766 3bit_freq_divider_1.sg13g2_tiehi_1.L_HI a_60584_24580# 0.12404f
C767 VDD a_53022_43738# 13.1862f
C768 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.nQ 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.Q 0.02712f
C769 3bit_freq_divider_1.freq_div_cell_0.Cin 3bit_freq_divider_1.sg13g2_tiehi_1.L_HI 0.14552f
C770 m4_17285_2698# Y0 0.3817f
C771 3bit_freq_divider_1.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 3bit_freq_divider_1.dff_nclk_0.D 0.17618f
C772 a_53065_20179# a_53445_20214# 0.41048f
C773 VDD a_52950_23913# 0.24052f
C774 VDD a_53899_24000# 0.26493f
C775 3bit_freq_divider_0.dff_nclk_0.nCLK a_53774_23690# 0.35198f
C776 m2_16847_2260# m1_16847_2260# 0.2063p
C777 3bit_freq_divider_0.dff_nclk_0.nCLK a_54504_23771# 0.37259f
C778 3bit_freq_divider_1.sg13g2_or3_1_0.C 3bit_freq_divider_1.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.28129f
C779 a_61887_24046# a_61691_24046# 0.45047f
C780 X0 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.Q 0.24362f
C781 VDD a_55770_40850# 0.01475f
C782 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.D 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.40308f
C783 X0 3bit_freq_divider_0.dff_nclk_0.D 0.1238f
C784 a_52950_23913# 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.nQ 0.21609f
C785 a_53065_23691# a_53774_23690# 0.02335f
C786 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.Q X1 0.15458f
C787 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.D a_61394_21976# 0.3562f
C788 VDD a_55769_40283# 1.37334f
C789 VDD m6_60810_42209# 0.03757f
C790 a_55862_56737# charge_pump_0.bias_p 0.3307f
C791 VDD 3bit_freq_divider_0.sg13g2_tiehi_1.L_HI 0.77158f
C792 VDD 3bit_freq_divider_1.dff_nclk_0.D 0.84615f
C793 a_62900_23691# VDD 0.31029f
C794 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 3bit_freq_divider_1.sg13g2_nand2_1_0.Y 0.11142f
C795 a_55969_42591# vco_wob_0.vctl 0.0811f
C796 X0 PFD_0.VCO_CLK 0.1115f
C797 VDD a_61394_20220# 0.36995f
C798 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.nQ a_53445_21970# 0.10118f
C799 VDD a_63255_21488# 0.26051f
C800 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.D 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.40308f
C801 a_52924_24641# 3bit_freq_divider_0.sg13g2_or3_1_0.C 0.10662f
C802 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.Q 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.D 0.22983f
C803 3bit_freq_divider_1.sg13g2_or3_1_0.C VDD 0.19202f
C804 Y2 a_63426_21130# 0.02209f
C805 a_51684_22692# VDD 0.19308f
C806 a_51648_24041# a_51631_22774# 0.02302f
C807 a_64383_23628# 3bit_freq_divider_1.dff_nclk_0.D 0.03728f
C808 m4_17285_2698# X0 0.39515f
C809 3bit_freq_divider_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK X1 0.02018f
C810 a_63426_24642# 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.Q 0.02246f
C811 a_53065_20179# a_53774_20178# 0.02335f
C812 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.Q a_54472_21129# 0.02559f
C813 VDD a_64384_21091# 0.34084f
C814 m5_17331_2744# CLK_OUT 0.40842f
C815 a_54494_43159# a_53022_43738# 0.04f
C816 X1 a_51693_23426# 0.01735f
C817 a_51684_22284# a_51684_22692# 0.47248f
C818 3bit_freq_divider_0.EN a_59097_54704# 0.03561f
C819 a_61707_23244# a_61878_22886# 0.36535f
C820 3bit_freq_divider_1.dff_nclk_0.nRST a_64731_24890# 0.01267f
C821 a_54627_42591# a_53152_43159# 0.03153f
C822 a_53065_21935# 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.Q 0.0119f
C823 a_54489_40413# a_53085_40283# 0.01232f
C824 3bit_freq_divider_1.freq_div_cell_0.Cout a_60967_21478# 0.13034f
C825 a_55345_23141# 3bit_freq_divider_0.freq_div_cell_0.Cout 0.13167f
C826 a_61878_22886# 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.Q 0.02559f
C827 3bit_freq_divider_1.freq_div_cell_0.Cout a_61707_21488# 0.12082f
C828 a_61394_21976# a_61887_22290# 0.47248f
C829 a_62270_20543# a_62654_20215# 0.03957f
C830 a_64383_23434# 3bit_freq_divider_1.dff_nclk_0.nRST 0.126f
C831 a_61394_23732# 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.D 0.3562f
C832 a_59097_54704# charge_pump_0.bias_p 0.04726f
C833 a_55345_24897# 3bit_freq_divider_0.sg13g2_tiehi_1.L_HI 0.21784f
C834 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.D 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.40308f
C835 a_62270_24055# 3bit_freq_divider_1.dff_nclk_0.nCLK 0.17312f
C836 a_64384_24445# CLK_OUT 0.1244f
C837 a_53065_21935# 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.nQ 0.0571f
C838 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.Q 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.nQ 0.02712f
C839 VDD 3bit_freq_divider_1.freq_div_cell_1.Cout 0.4595f
C840 3bit_freq_divider_1.dff_nclk_0.nCLK a_62654_20215# 0.31114f
C841 a_64383_23706# 3bit_freq_divider_1.dff_nclk_0.D 0.12409f
C842 a_53738_20514# a_53899_20488# 0.66077f
C843 a_52886_23148# 3bit_freq_divider_0.sg13g2_or3_1_0.B 0.23215f
C844 X0 m1_17285_2698# 0.01061f
C845 3bit_freq_divider_0.EN nEN 0.24728f
C846 Y2 a_62654_23727# 0.02178f
C847 a_56695_49467# charge_pump_0.vout 0.02916f
C848 3bit_freq_divider_0.freq_div_cell_1.Cout a_54434_21392# 0.01154f
C849 3bit_freq_divider_0.EN 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.D 0.02119f
C850 3bit_freq_divider_0.freq_div_cell_0.Cout VDD 1.22849f
C851 a_63255_25000# Y2 0.02709f
C852 3bit_freq_divider_1.dff_nclk_0.nCLK 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.nQ 0.02503f
C853 Y2 a_63463_21972# 0.01788f
C854 3bit_freq_divider_1.sg13g2_or3_1_0.B 3bit_freq_divider_1.sg13g2_or3_1_0.A 0.72102f
C855 CLK_IN m3_17285_2698# 0.30224f
C856 a_61878_24642# 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.Q 0.02559f
C857 a_53147_40413# a_54428_40850# 0.23834f
C858 a_51648_24438# 3bit_freq_divider_0.dff_nclk_0.D 0.2233f
C859 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.nQ Y1 0.01108f
C860 nEN charge_pump_0.bias_p 0.0229f
C861 a_53350_24641# a_52886_24904# 0.0104f
C862 vco_wob_0.vctl a_53086_40850# 0.04284f
C863 3bit_freq_divider_1.dff_nclk_0.nCLK a_63463_20216# 0.05882f
C864 a_58536_54976# charge_pump_0.bias_n 0.02549f
C865 3bit_freq_divider_0.dff_nclk_0.nCLK a_53065_20179# 0.31132f
C866 a_51684_22692# 3bit_freq_divider_0.dff_nclk_0.nRST 0.126f
C867 a_54427_40283# a_53147_40413# 0.42019f
C868 3bit_freq_divider_0.sg13g2_or3_1_0.B 3bit_freq_divider_0.dff_nclk_0.nCLK 0.58488f
C869 Y2 a_63255_23244# 0.01433f
C870 a_62119_22361# a_61394_21976# 0.45825f
C871 a_54472_22885# a_54434_23148# 0.36535f
C872 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.D 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.Q 0.22983f
C873 a_46817_27899# a_47954_28913# 0.22374f
C874 a_51648_24438# PFD_0.VCO_CLK 0.11636f
C875 a_55969_42591# VDD 0.0108f
C876 VDD a_61887_20534# 0.19386f
C877 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.sg13g2_dfrbp_1_0.CLK a_53738_20514# 0.01324f
C878 a_55862_56737# VDD 0.47223f
C879 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 3bit_freq_divider_0.sg13g2_nand2_1_0.Y 0.10521f
C880 3bit_freq_divider_1.sg13g2_or3_1_0.C a_63426_24642# 0.10662f
C881 3bit_freq_divider_1.dff_nclk_0.nCLK 3bit_freq_divider_1.freq_div_cell_0.Cout 0.32366f
C882 3bit_freq_divider_1.sg13g2_nand2_1_0.Y 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.10521f
C883 a_60528_49446# vco_wob_0.vctl 0.01545f
C884 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.D a_61394_20220# 0.3562f
C885 VDD a_51708_21299# 0.01263f
C886 a_64362_24865# a_64731_24890# 0.01952f
C887 m2_17285_2698# m3_17285_2698# 0.20496p
C888 a_53968_23946# a_53774_23690# 0.05314f
C889 a_53968_23946# a_54504_23771# 0.45825f
C890 3bit_freq_divider_1.freq_div_cell_0.Cin 3bit_freq_divider_1.freq_div_cell_0.Cout 0.10559f
C891 a_58454_40850# a_58515_40413# 0.03243f
C892 a_61878_24642# 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.D 0.12185f
C893 m7_16847_2260# CLK_OUT 1.40976f
C894 m4_17285_2698# Y1 0.3817f
C895 3bit_freq_divider_0.freq_div_cell_1.Cout 3bit_freq_divider_0.sg13g2_nand2_1_0.Y 0.07626f
C896 VDD a_60385_24947# 0.11858f
C897 a_64383_23434# 3bit_freq_divider_1.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.01473f
C898 a_57178_43159# vco_wob_0.vctl 0.026f
C899 a_51685_23725# 3bit_freq_divider_0.dff_nclk_0.D 0.12409f
C900 a_64419_23326# a_64383_23300# 0.70262f
C901 a_56887_49467# charge_pump_0.vout 0.63953f
C902 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.Q X1 0.01869f
C903 3bit_freq_divider_0.EN charge_pump_0.bias_p 0.33628f
C904 a_53738_22270# a_54504_22015# 0.47248f
C905 a_61887_24046# a_62900_23691# 0.04306f
C906 Y0 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.Q 0.20944f
C907 a_53774_21934# a_53738_22270# 0.44698f
C908 a_52944_43077# a_53022_43738# 0.93638f
C909 3bit_freq_divider_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 3bit_freq_divider_0.sg13g2_or3_1_0.C 0.28129f
C910 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.D 3bit_freq_divider_1.freq_div_cell_0.Cout 0.084f
C911 VDD a_64731_24890# 0.04155f
C912 VDD a_53085_40283# 1.35573f
C913 3bit_freq_divider_0.dff_nclk_0.D X1 0.11556f
C914 a_61707_23244# 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.Q 0.46099f
C915 VDD a_63426_21130# 0.20953f
C916 a_61691_20534# a_62654_20215# 0.02302f
C917 3bit_freq_divider_0.dff_nclk_0.nCLK a_52950_20401# 0.05883f
C918 VDD 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.30706f
C919 a_64383_23434# VDD 0.19308f
C920 PFD_0.DOWN PFD_0.UP 0.20773f
C921 3bit_freq_divider_0.EN X2 0.11756f
C922 a_55969_42591# a_54494_43159# 0.03153f
C923 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.D VDD 0.97078f
C924 VDD a_59799_40285# 1.38295f
C925 3bit_freq_divider_1.freq_div_cell_1.Cout 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.D 0.04623f
C926 a_63463_23728# 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.nQ 0.21609f
C927 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.D 3bit_freq_divider_1.sg13g2_nand2_1_0.Y 0.04726f
C928 3bit_freq_divider_1.dff_nclk_0.nCLK 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.60301f
C929 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 3bit_freq_divider_0.sg13g2_nand2_1_0.Y 0.11142f
C930 a_52944_43077# a_53285_42591# 0.03491f
C931 VDD a_61707_25000# 0.27566f
C932 a_60385_24717# a_60385_24947# 0.10864f
C933 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.D 3bit_freq_divider_0.sg13g2_nand2_1_0.Y 0.05125f
C934 3bit_freq_divider_1.dff_nclk_0.nCLK 3bit_freq_divider_1.sg13g2_or3_1_0.A 0.48568f
C935 3bit_freq_divider_1.dff_nclk_0.D a_64384_24445# 0.2233f
C936 a_54489_40413# vco_wob_0.vctl 0.04184f
C937 a_53022_43738# a_53058_43159# 0.24146f
C938 a_64383_23434# a_64383_23628# 0.44985f
C939 3bit_freq_divider_0.dff_nclk_0.nCLK a_53899_24000# 0.17312f
C940 a_57084_43159# a_53022_43738# 0.19696f
C941 VDD a_53968_20434# 0.2982f
C942 3bit_freq_divider_0.EN CLK_IN 0.09396f
C943 a_51684_22692# a_51648_24041# 0.40027f
C944 a_53774_21934# a_54504_22015# 0.17766f
C945 nEN VDD 3.87548f
C946 PFD_0.DOWN PFD_0.VCO_CLK 0.20401f
C947 a_52950_23913# a_53065_23691# 0.09575f
C948 a_53065_23691# a_53899_24000# 0.03957f
C949 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.D 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.40308f
C950 VDD a_60967_24990# 0.4548f
C951 VDD 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.D 0.9437f
C952 X0 a_52886_24904# 0.40762f
C953 a_64424_22200# a_64383_23300# 0.45825f
C954 a_62654_21971# 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.nQ 0.0571f
C955 a_62654_23727# VDD 0.43765f
C956 a_57111_40283# a_53022_43738# 0.18962f
C957 charge_pump_0.bias_p a_54357_49278# 0.01013f
C958 3bit_freq_divider_1.dff_nclk_0.nCLK a_61691_24046# 0.35198f
C959 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.Q a_60967_21478# 0.30546f
C960 a_58653_42591# 3bit_freq_divider_0.CLK_IN 0.2448f
C961 a_59800_40852# vco_wob_0.vctl 0.05123f
C962 a_58536_54976# a_58734_56203# 0.19076f
C963 3bit_freq_divider_1.freq_div_cell_0.Cout a_61878_21130# 0.01011f
C964 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.Q a_62654_21971# 0.0119f
C965 a_63255_25000# VDD 0.26507f
C966 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.Q a_61707_21488# 0.46099f
C967 VDD a_63463_21972# 0.2345f
C968 a_55862_56737# a_55948_56737# 0.0609f
C969 a_64383_23434# a_64383_23706# 0.04306f
C970 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.Q 3bit_freq_divider_0.CLK_IN 0.02001f
C971 3bit_freq_divider_1.sg13g2_or3_1_0.C Y0 0.12518f
C972 CLK_IN a_46749_30782# 0.97391f
C973 VDD a_57178_43159# 1.11494f
C974 a_63255_23244# VDD 0.25835f
C975 a_53738_22270# VDD 0.21577f
C976 3bit_freq_divider_1.dff_nclk_0.nCLK a_62900_20179# 0.2629f
C977 a_47777_29803# PFD_0.UP 0.62819f
C978 3bit_freq_divider_1.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 3bit_freq_divider_1.dff_nclk_0.nRST 0.16234f
C979 a_51693_23075# VDD 0.2446f
C980 Y2 VDD 1.18034f
C981 a_45658_27900# PFD_0.DOWN 0.61911f
C982 3bit_freq_divider_1.dff_nclk_0.nRST a_64362_24865# 0.03098f
C983 a_55345_21385# VDD 0.45855f
C984 X2 3bit_freq_divider_0.sg13g2_or3_1_0.A 0.2051f
C985 3bit_freq_divider_0.EN VDD 6.40652f
C986 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.Q 3bit_freq_divider_0.freq_div_cell_0.Cin 0.42266f
C987 a_58426_43159# 3bit_freq_divider_0.CLK_IN 0.4131f
C988 a_57173_40413# vco_wob_0.vctl 0.03129f
C989 a_62270_20543# a_62119_20605# 0.70262f
C990 a_52924_24641# 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.Q 0.02246f
C991 CLK_IN m6_17427_2840# 1.23795f
C992 CLK_OUT Y1 0.01478f
C993 a_51685_23725# a_51631_22774# 0.04324f
C994 a_61887_22290# 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.01324f
C995 3bit_freq_divider_0.sg13g2_or3_1_0.C a_51648_21103# 0.25034f
C996 a_56013_24979# 3bit_freq_divider_0.sg13g2_tiehi_1.L_HI 0.02161f
C997 3bit_freq_divider_0.sg13g2_or3_1_0.C 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.Q 0.05745f
C998 VDD a_62270_22299# 0.26052f
C999 3bit_freq_divider_1.dff_nclk_0.nCLK 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.nQ 0.0874f
C1000 3bit_freq_divider_1.sg13g2_nand2_1_0.Y 3bit_freq_divider_1.freq_div_cell_1.Cout 0.07626f
C1001 VDD charge_pump_0.bias_p 2.67087f
C1002 VDD 3bit_freq_divider_1.dff_nclk_0.nRST 0.60883f
C1003 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.Q a_53065_20179# 0.01984f
C1004 3bit_freq_divider_1.dff_nclk_0.nCLK a_62119_20605# 0.32732f
C1005 X1 a_51631_22774# 0.02271f
C1006 VDD a_54489_40413# 1.15543f
C1007 a_51708_21413# a_51648_21103# 0.014f
C1008 3bit_freq_divider_1.dff_nclk_0.nCLK 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.60301f
C1009 3bit_freq_divider_1.dff_nclk_0.nCLK 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.Q 1.04018f
C1010 a_60967_23234# VDD 0.45855f
C1011 VDD vco_wob_0.vctl 0.2823f
C1012 3bit_freq_divider_0.freq_div_cell_0.Cout 3bit_freq_divider_0.dff_nclk_0.nCLK 0.32366f
C1013 3bit_freq_divider_0.CLK_IN a_53022_43738# 0.16863f
C1014 a_54504_22015# VDD 0.38024f
C1015 a_53774_21934# VDD 0.69275f
C1016 3bit_freq_divider_1.sg13g2_or3_1_0.C 3bit_freq_divider_1.sg13g2_or3_1_0.B 1.00414f
C1017 m5_16847_2260# m4_16847_2260# 0.2063p
C1018 VDD a_46749_30782# 1.12191f
C1019 a_51759_25014# a_51721_24988# 0.10864f
C1020 a_64383_23628# 3bit_freq_divider_1.dff_nclk_0.nRST 0.3268f
C1021 X2 VDD 0.25402f
C1022 3bit_freq_divider_1.dff_nclk_0.nCLK 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.Q 0.0844f
C1023 a_54434_21392# a_54472_21129# 0.36535f
C1024 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.Q Y1 0.18013f
C1025 3bit_freq_divider_1.sg13g2_or3_1_0.B a_64384_21091# 0.26158f
C1026 a_62270_22299# a_61691_22290# 0.04304f
C1027 3bit_freq_divider_1.freq_div_cell_0.Cin 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.Q 0.22232f
C1028 a_53065_21935# 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.Q 0.01984f
C1029 a_53445_23726# VDD 0.31261f
C1030 a_62119_24117# VDD 0.32287f
C1031 a_63255_25000# a_63426_24642# 0.36535f
C1032 m6_60810_42209# 3bit_freq_divider_0.CLK_IN 0.11742f
C1033 3bit_freq_divider_0.sg13g2_or3_1_0.B X1 0.27832f
C1034 a_56695_49467# a_56887_49467# 0.01287f
C1035 3bit_freq_divider_0.freq_div_cell_0.Cin 3bit_freq_divider_0.sg13g2_nand2_1_0.Y 0.25573f
C1036 a_51693_23075# 3bit_freq_divider_0.dff_nclk_0.nRST 0.16442f
C1037 CLK_IN VDD 2.49441f
C1038 VDD a_54357_49278# 0.31963f
C1039 m2_16847_2260# m3_16847_2260# 0.2063p
C1040 a_53774_20178# a_53968_20434# 0.05314f
C1041 a_53065_20179# a_53899_20488# 0.03957f
C1042 a_53968_23946# a_53899_24000# 0.70262f
C1043 a_53445_23726# 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.nQ 0.10118f
C1044 a_53738_24026# a_53774_23690# 0.44698f
C1045 a_53738_24026# a_54504_23771# 0.47248f
C1046 a_53085_40283# a_52944_43077# 0.45412f
C1047 a_62900_20179# a_61691_20534# 0.04324f
C1048 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.Q a_52950_20401# 0.12389f
C1049 a_61878_24642# a_61707_25000# 0.36535f
C1050 a_55941_24882# 3bit_freq_divider_0.sg13g2_tiehi_1.L_HI 0.12404f
C1051 3bit_freq_divider_1.dff_nclk_0.nCLK 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.D 0.21603f
C1052 VDD 3bit_freq_divider_0.sg13g2_or3_1_0.A 0.12791f
C1053 3bit_freq_divider_0.freq_div_cell_0.Cout a_54434_23148# 0.01154f
C1054 a_64383_23706# 3bit_freq_divider_1.dff_nclk_0.nRST 0.25925f
C1055 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.D a_53774_20178# 0.01446f
C1056 a_54494_43159# vco_wob_0.vctl 0.0248f
C1057 a_61887_24046# a_62654_23727# 0.40027f
C1058 3bit_freq_divider_1.freq_div_cell_0.Cin 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.D 0.084f
C1059 a_53065_21935# a_53445_21970# 0.41048f
C1060 a_55345_23141# VDD 0.45855f
C1061 3bit_freq_divider_1.dff_nclk_0.sg13g2_dfrbp_1_0.CLK VDD 0.28742f
C1062 VDD a_64362_24865# 0.08341f
C1063 a_61707_23244# 3bit_freq_divider_1.freq_div_cell_0.Cout 0.01154f
C1064 3bit_freq_divider_0.EN 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.D 0.02092f
C1065 VDD a_57173_40413# 0.98193f
C1066 a_45579_29803# a_45451_28860# 0.44406f
C1067 3bit_freq_divider_1.freq_div_cell_0.Cout 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.Q 0.22232f
C1068 a_61691_20534# a_62119_20605# 0.05314f
C1069 Y0 m3_17285_2698# 0.2919f
C1070 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.nQ a_62900_21935# 0.10118f
C1071 3bit_freq_divider_0.EN a_55948_56737# 0.0294f
C1072 3bit_freq_divider_0.dff_nclk_0.nCLK 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.sg13g2_dfrbp_1_0.CLK 0.60301f
C1073 a_56742_53480# a_56828_53480# 0.09853f
C1074 VDD 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.nQ 0.18065f
C1075 a_60967_21478# 3bit_freq_divider_1.freq_div_cell_1.Cout 0.13166f
C1076 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.sg13g2_dfrbp_1_0.CLK a_61691_20534# 0.33731f
C1077 3bit_freq_divider_1.dff_nclk_0.sg13g2_dfrbp_1_0.CLK a_64383_23628# 0.33833f
C1078 3bit_freq_divider_1.dff_nclk_0.nCLK 3bit_freq_divider_1.dff_nclk_0.D 0.04354f
C1079 3bit_freq_divider_0.dff_nclk_0.nCLK 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.D 0.21603f
C1080 3bit_freq_divider_1.freq_div_cell_1.Cout a_61707_21488# 0.01154f
C1081 a_52944_43077# a_53086_40850# 0.23665f
C1082 3bit_freq_divider_1.dff_nclk_0.nCLK a_62900_23691# 0.24211f
C1083 Y2 VSS 0.12039p
C1084 X2 VSS 91.68561f
C1085 Y1 VSS 0.10102p
C1086 X1 VSS 94.7177f
C1087 CLK_OUT VSS 92.2343f
C1088 Y0 VSS 92.142f
C1089 X0 VSS 90.2415f
C1090 CLK_IN VSS 93.6639f
C1091 nEN VSS 0.10244p
C1092 VDD VSS 0.19687p
C1093 m7_16847_2260# VSS 93.0612f
C1094 m6_60810_42209# VSS 1.80367f
C1095 m6_17427_2840# VSS 0.10708p
C1096 m6_16847_2260# VSS 0.11472p
C1097 m5_17331_2744# VSS 79.2024f
C1098 m5_16847_2260# VSS 84.4749f
C1099 m4_17285_2698# VSS 84.41901f
C1100 m4_16847_2260# VSS 89.24989f
C1101 m3_17285_2698# VSS 91.8291f
C1102 m3_16847_2260# VSS 96.21301f
C1103 m2_17285_2698# VSS 0.10557p
C1104 m2_16847_2260# VSS 0.10679p
C1105 m1_17285_2698# VSS 0.22685p
C1106 m1_16847_2260# VSS 0.22893p
C1107 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.nQ VSS 0.08893f $ **FLOATING
C1108 a_62900_20179# VSS 0.34783f $ **FLOATING
C1109 a_63463_20216# VSS 0.43565f $ **FLOATING
C1110 a_62654_20215# VSS 0.80634f $ **FLOATING
C1111 a_62119_20605# VSS 0.26895f $ **FLOATING
C1112 a_62270_20543# VSS 0.16883f $ **FLOATING
C1113 a_61887_20534# VSS 1.05953f $ **FLOATING
C1114 a_61394_20220# VSS 0.13262f $ **FLOATING
C1115 a_61691_20534# VSS 0.79964f $ **FLOATING
C1116 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.sg13g2_dfrbp_1_0.CLK VSS 0.51487f $ **FLOATING
C1117 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.sg13g2_dfrbp_1_0.CLK VSS 0.51489f $ **FLOATING
C1118 a_54504_20259# VSS 0.13262f $ **FLOATING
C1119 a_53899_20488# VSS 0.16883f $ **FLOATING
C1120 a_53968_20434# VSS 0.26896f $ **FLOATING
C1121 a_53738_20514# VSS 1.05953f $ **FLOATING
C1122 a_53445_20214# VSS 0.34783f $ **FLOATING
C1123 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.nQ VSS 0.08893f $ **FLOATING
C1124 a_53774_20178# VSS 0.80054f $ **FLOATING
C1125 a_53065_20179# VSS 0.80634f $ **FLOATING
C1126 a_52950_20401# VSS 0.43566f $ **FLOATING
C1127 a_64384_21091# VSS 0.59054f $ **FLOATING
C1128 3bit_freq_divider_1.sg13g2_or3_1_0.A VSS 0.77543f $ **FLOATING
C1129 a_63255_21488# VSS 0.38381f $ **FLOATING
C1130 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.D VSS 0.49782f $ **FLOATING
C1131 a_61707_21488# VSS 0.36496f $ **FLOATING
C1132 3bit_freq_divider_1.freq_div_cell_1.Cout VSS 0.14556f $ **FLOATING
C1133 a_60967_21478# VSS 0.27989f $ **FLOATING
C1134 3bit_freq_divider_1.freq_div_cell_1.dff_nclk_0.Q VSS 2.25165f $ **FLOATING
C1135 3bit_freq_divider_0.freq_div_cell_1.Cout VSS 0.14556f $ **FLOATING
C1136 a_55345_21385# VSS 0.27989f $ **FLOATING
C1137 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.D VSS 0.49784f $ **FLOATING
C1138 a_54434_21392# VSS 0.36496f $ **FLOATING
C1139 3bit_freq_divider_0.sg13g2_or3_1_0.A VSS 0.77447f $ **FLOATING
C1140 a_51648_21103# VSS 0.59026f $ **FLOATING
C1141 a_52886_21392# VSS 0.3838f $ **FLOATING
C1142 3bit_freq_divider_0.freq_div_cell_1.dff_nclk_0.Q VSS 2.25169f $ **FLOATING
C1143 a_60922_21796# VSS 0.03012f $ **FLOATING
C1144 a_60922_21818# VSS 0.02768f $ **FLOATING
C1145 a_52808_21795# VSS 0.03012f $ **FLOATING
C1146 a_52808_21817# VSS 0.02768f $ **FLOATING
C1147 3bit_freq_divider_1.dff_nclk_0.sg13g2_dfrbp_1_0.CLK VSS 0.50854f $ **FLOATING
C1148 a_64424_22200# VSS 0.12168f $ **FLOATING
C1149 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.nQ VSS 0.07921f $ **FLOATING
C1150 a_62900_21935# VSS 0.33549f $ **FLOATING
C1151 a_63463_21972# VSS 0.42316f $ **FLOATING
C1152 a_62654_21971# VSS 0.7639f $ **FLOATING
C1153 a_62119_22361# VSS 0.25006f $ **FLOATING
C1154 a_62270_22299# VSS 0.1501f $ **FLOATING
C1155 a_61887_22290# VSS 1.02135f $ **FLOATING
C1156 a_61394_21976# VSS 0.12168f $ **FLOATING
C1157 a_61691_22290# VSS 0.77938f $ **FLOATING
C1158 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK VSS 0.47143f $ **FLOATING
C1159 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK VSS 0.47143f $ **FLOATING
C1160 a_54504_22015# VSS 0.12168f $ **FLOATING
C1161 a_53899_22244# VSS 0.1501f $ **FLOATING
C1162 a_53968_22190# VSS 0.25006f $ **FLOATING
C1163 a_53738_22270# VSS 1.02135f $ **FLOATING
C1164 a_53445_21970# VSS 0.33549f $ **FLOATING
C1165 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.nQ VSS 0.07921f $ **FLOATING
C1166 a_53774_21934# VSS 0.78026f $ **FLOATING
C1167 a_53065_21935# VSS 0.7639f $ **FLOATING
C1168 a_52950_22157# VSS 0.4233f $ **FLOATING
C1169 3bit_freq_divider_1.sg13g2_or3_1_0.B VSS 1.39257f $ **FLOATING
C1170 a_64383_23300# VSS 0.25093f $ **FLOATING
C1171 a_63255_23244# VSS 0.37914f $ **FLOATING
C1172 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.D VSS 0.45601f $ **FLOATING
C1173 a_61707_23244# VSS 0.36159f $ **FLOATING
C1174 3bit_freq_divider_1.freq_div_cell_0.Cout VSS 1.80113f $ **FLOATING
C1175 a_60967_23234# VSS 0.27786f $ **FLOATING
C1176 a_64419_23326# VSS 0.1501f $ **FLOATING
C1177 3bit_freq_divider_1.freq_div_cell_0.dff_nclk_0.Q VSS 2.24178f $ **FLOATING
C1178 3bit_freq_divider_0.dff_nclk_0.sg13g2_dfrbp_1_0.CLK VSS 0.50854f $ **FLOATING
C1179 a_51684_22284# VSS 0.12168f $ **FLOATING
C1180 3bit_freq_divider_0.freq_div_cell_0.Cout VSS 1.80115f $ **FLOATING
C1181 a_55345_23141# VSS 0.27786f $ **FLOATING
C1182 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.D VSS 0.45601f $ **FLOATING
C1183 a_54434_23148# VSS 0.36159f $ **FLOATING
C1184 3bit_freq_divider_0.sg13g2_or3_1_0.B VSS 1.39146f $ **FLOATING
C1185 a_52886_23148# VSS 0.37912f $ **FLOATING
C1186 3bit_freq_divider_0.freq_div_cell_0.dff_nclk_0.Q VSS 2.2418f $ **FLOATING
C1187 a_64383_23628# VSS 0.82074f $ **FLOATING
C1188 a_64383_23434# VSS 1.02665f $ **FLOATING
C1189 a_60922_23552# VSS 0.03012f $ **FLOATING
C1190 a_60922_23574# VSS 0.02768f $ **FLOATING
C1191 a_52808_23551# VSS 0.03012f $ **FLOATING
C1192 a_52808_23573# VSS 0.02768f $ **FLOATING
C1193 a_51693_23426# VSS 0.25093f $ **FLOATING
C1194 a_51693_23075# VSS 0.1501f $ **FLOATING
C1195 a_64383_23706# VSS 0.33666f $ **FLOATING
C1196 3bit_freq_divider_1.dff_nclk_0.D VSS 0.57206f $ **FLOATING
C1197 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.nQ VSS 0.08281f $ **FLOATING
C1198 a_62900_23691# VSS 0.33612f $ **FLOATING
C1199 a_63463_23728# VSS 0.42235f $ **FLOATING
C1200 a_62654_23727# VSS 0.76426f $ **FLOATING
C1201 a_62119_24117# VSS 0.25006f $ **FLOATING
C1202 a_62270_24055# VSS 0.1501f $ **FLOATING
C1203 a_61887_24046# VSS 1.02191f $ **FLOATING
C1204 a_61394_23732# VSS 0.12168f $ **FLOATING
C1205 a_61691_24046# VSS 0.78738f $ **FLOATING
C1206 3bit_freq_divider_1.dff_nclk_0.nCLK VSS 7.48134f $ **FLOATING
C1207 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.sg13g2_dfrbp_1_0.CLK VSS 0.47246f $ **FLOATING
C1208 a_51631_22774# VSS 0.82147f $ **FLOATING
C1209 a_51684_22692# VSS 1.02713f $ **FLOATING
C1210 3bit_freq_divider_1.sg13g2_nand2_1_0.Y VSS 2.56526f $ **FLOATING
C1211 3bit_freq_divider_0.sg13g2_nand2_1_0.Y VSS 2.56527f $ **FLOATING
C1212 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.sg13g2_dfrbp_1_0.CLK VSS 0.47246f $ **FLOATING
C1213 a_54504_23771# VSS 0.12168f $ **FLOATING
C1214 a_53899_24000# VSS 0.1501f $ **FLOATING
C1215 a_53968_23946# VSS 0.25006f $ **FLOATING
C1216 a_53738_24026# VSS 1.02191f $ **FLOATING
C1217 a_53445_23726# VSS 0.33612f $ **FLOATING
C1218 3bit_freq_divider_0.dff_nclk_0.nCLK VSS 7.50548f $ **FLOATING
C1219 a_51685_23725# VSS 0.33666f $ **FLOATING
C1220 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.nQ VSS 0.08281f $ **FLOATING
C1221 a_53774_23690# VSS 0.78853f $ **FLOATING
C1222 a_53065_23691# VSS 0.76426f $ **FLOATING
C1223 a_52950_23913# VSS 0.42231f $ **FLOATING
C1224 a_64383_23889# VSS 0.79267f $ **FLOATING
C1225 a_64384_24445# VSS 0.41218f $ **FLOATING
C1226 3bit_freq_divider_0.dff_nclk_0.D VSS 0.57206f $ **FLOATING
C1227 a_51648_24041# VSS 0.7928f $ **FLOATING
C1228 3bit_freq_divider_1.dff_nclk_0.nRST VSS 1.21235f $ **FLOATING
C1229 a_64398_24796# VSS 0.17085f $ **FLOATING
C1230 a_64338_24910# VSS 0.01158f $ **FLOATING
C1231 a_64362_24865# VSS 0.18902f $ **FLOATING
C1232 a_64459_24995# VSS 0.21807f $ **FLOATING
C1233 a_51648_24438# VSS 0.41218f $ **FLOATING
C1234 3bit_freq_divider_1.sg13g2_or3_1_0.C VSS 2.00849f $ **FLOATING
C1235 a_63255_25000# VSS 0.38174f $ **FLOATING
C1236 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.D VSS 0.4595f $ **FLOATING
C1237 a_61707_25000# VSS 0.36409f $ **FLOATING
C1238 3bit_freq_divider_1.freq_div_cell_0.Cin VSS 1.81006f $ **FLOATING
C1239 a_60967_24990# VSS 0.27856f $ **FLOATING
C1240 3bit_freq_divider_1.freq_div_cell_2.dff_nclk_0.Q VSS 2.27033f $ **FLOATING
C1241 a_60584_24580# VSS 0.16608f $ **FLOATING
C1242 a_60385_24947# VSS 0.21087f $ **FLOATING
C1243 a_56137_24678# VSS 0.21087f $ **FLOATING
C1244 3bit_freq_divider_1.sg13g2_tiehi_1.L_HI VSS 1.60229f $ **FLOATING
C1245 a_60385_24717# VSS 0.17977f $ **FLOATING
C1246 a_60479_25023# VSS 0.01118f $ **FLOATING
C1247 a_55941_24882# VSS 0.16608f $ **FLOATING
C1248 3bit_freq_divider_0.dff_nclk_0.nRST VSS 1.20799f $ **FLOATING
C1249 a_51622_24863# VSS 0.17085f $ **FLOATING
C1250 3bit_freq_divider_0.freq_div_cell_0.Cin VSS 1.81006f $ **FLOATING
C1251 a_55345_24897# VSS 0.27856f $ **FLOATING
C1252 a_56039_25022# VSS 0.01118f $ **FLOATING
C1253 a_56013_24979# VSS 0.17977f $ **FLOATING
C1254 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.D VSS 0.4595f $ **FLOATING
C1255 a_54434_24904# VSS 0.36409f $ **FLOATING
C1256 3bit_freq_divider_0.sg13g2_or3_1_0.C VSS 2.00844f $ **FLOATING
C1257 a_52065_24890# VSS 0.01158f $ **FLOATING
C1258 a_51721_24988# VSS 0.21807f $ **FLOATING
C1259 a_51759_25014# VSS 0.18902f $ **FLOATING
C1260 a_52886_24904# VSS 0.38144f $ **FLOATING
C1261 3bit_freq_divider_0.sg13g2_tiehi_1.L_HI VSS 1.60229f $ **FLOATING
C1262 3bit_freq_divider_0.freq_div_cell_2.dff_nclk_0.Q VSS 2.27033f $ **FLOATING
C1263 a_47954_28913# VSS 0.97627f $ **FLOATING
C1264 a_46817_27899# VSS 1.26528f $ **FLOATING
C1265 a_45658_27900# VSS 1.24513f $ **FLOATING
C1266 PFD_0.VCO_CLK VSS 5.09845f $ **FLOATING
C1267 a_48909_28913# VSS 1.03223f $ **FLOATING
C1268 a_45451_28860# VSS 1.00878f $ **FLOATING
C1269 a_47777_29803# VSS 1.2524f $ **FLOATING
C1270 a_46749_30782# VSS 1.31435f $ **FLOATING
C1271 a_45579_29803# VSS 0.97532f $ **FLOATING
C1272 a_59799_40285# VSS 0.05072f $ **FLOATING
C1273 a_58453_40283# VSS 0.04654f $ **FLOATING
C1274 a_57111_40283# VSS 0.0474f $ **FLOATING
C1275 a_55769_40283# VSS 0.04814f $ **FLOATING
C1276 a_54427_40283# VSS 0.04567f $ **FLOATING
C1277 a_53085_40283# VSS 0.07408f $ **FLOATING
C1278 a_58515_40413# VSS 4.51596f $ **FLOATING
C1279 a_57173_40413# VSS 4.66235f $ **FLOATING
C1280 a_55831_40413# VSS 4.71205f $ **FLOATING
C1281 a_54489_40413# VSS 5.15226f $ **FLOATING
C1282 a_53147_40413# VSS 5.26745f $ **FLOATING
C1283 a_59800_40852# VSS 0.75306f $ **FLOATING
C1284 a_58454_40850# VSS 0.8045f $ **FLOATING
C1285 a_57112_40850# VSS 0.81785f $ **FLOATING
C1286 a_55770_40850# VSS 0.82955f $ **FLOATING
C1287 a_54428_40850# VSS 0.82862f $ **FLOATING
C1288 a_53086_40850# VSS 0.83893f $ **FLOATING
C1289 a_58653_42591# VSS 0.65187f $ **FLOATING
C1290 a_57311_42591# VSS 0.67139f $ **FLOATING
C1291 a_55969_42591# VSS 0.6715f $ **FLOATING
C1292 a_54627_42591# VSS 0.67644f $ **FLOATING
C1293 a_53285_42591# VSS 0.68389f $ **FLOATING
C1294 3bit_freq_divider_0.CLK_IN VSS 20.6212f $ **FLOATING
C1295 a_57178_43159# VSS 5.00808f $ **FLOATING
C1296 a_55836_43159# VSS 4.39926f $ **FLOATING
C1297 a_54494_43159# VSS 4.398f $ **FLOATING
C1298 a_53152_43159# VSS 4.66518f $ **FLOATING
C1299 a_52944_43077# VSS 6.1695f $ **FLOATING
C1300 a_58426_43159# VSS 0.05888f $ **FLOATING
C1301 a_57084_43159# VSS 0.03844f $ **FLOATING
C1302 a_55742_43159# VSS 0.04051f $ **FLOATING
C1303 a_54400_43159# VSS 0.04084f $ **FLOATING
C1304 a_53058_43159# VSS 0.05472f $ **FLOATING
C1305 a_53022_43738# VSS 5.68098f $ **FLOATING
C1306 a_54747_49259# VSS 0.16684f $ **FLOATING
C1307 PFD_0.DOWN VSS 13.9137f $ **FLOATING
C1308 a_60528_49446# VSS 0.16044f
C1309 a_56695_49467# VSS 0.14015f
C1310 vco_wob_0.vctl VSS 17.2852f $ **FLOATING
C1311 a_56887_49467# VSS 8.04158f $ **FLOATING
C1312 a_54357_49278# VSS 0.26592f $ **FLOATING
C1313 PFD_0.UP VSS 12.6721f $ **FLOATING
C1314 charge_pump_0.vout VSS 28.7608f $ **FLOATING
C1315 a_56828_53480# VSS 2.32258f
C1316 a_56742_53480# VSS 1.67237f $ **FLOATING
C1317 a_59097_54704# VSS 0.1681f $ **FLOATING
C1318 a_58536_54976# VSS 0.61525f $ **FLOATING
C1319 a_58734_56203# VSS 0.05948f $ **FLOATING
C1320 charge_pump_0.bias_p VSS 5.47872f $ **FLOATING
C1321 charge_pump_0.bias_n VSS 6.55127f $ **FLOATING
C1322 3bit_freq_divider_0.EN VSS 51.6717f $ **FLOATING
C1323 a_55948_56737# VSS 1.95792f
C1324 a_55862_56737# VSS 0.99714f $ **FLOATING
.ends
