* Extracted by KLayout with SG13G2 LVS runset on : 02/09/2025 16:28

.SUBCKT FMD_QNC_PLL_3BIT_DIV
X$1 \$1 \$1 \$47 \$7 \$42 \$45 \$9 \$9 Bias_gen
X$24616 \$9 \$1 \$10 \$11 \$44 \$12 PFD
X$28388 \$1 \$43 \$28 loop_filter
X$29064 \$9 \$1 \$47 \$7 sg13g2_inv_1
X$33458 \$1 \$9 \$I71949 \$7 \$8 sg13g2_nand2_1
X$33459 \$9 \$1 \$I71956 sg13g2_tiehi
X$33460 \$11 \$I71954 \$I71954 \$I71950 \$1 \$I71956 \$9 dff_nclk
X$33461 \$1 \$9 \$I71950 \$I71951 \$I71953 \$I71952 sg13g2_or3_1
X$33462 \$I71951 \$2 \$I71949 \$I71955 \$I71958 \$1 \$I71950 \$9 freq_div_cell
X$33463 \$I71952 \$5 \$I71949 \$I71958 \$I71957 \$1 \$I71950 \$9 freq_div_cell
X$33464 \$9 \$1 \$I71957 sg13g2_tiehi
X$33465 \$I71953 \$3 \$I71949 \$I71959 \$I71955 \$1 \$I71950 \$9 freq_div_cell
X$33466 \$1 \$9 \$I71960 \$7 \$8 sg13g2_nand2_1
X$33467 \$9 \$1 \$I71967 sg13g2_tiehi
X$33468 \$6 \$I71965 \$I71965 \$I71961 \$1 \$I71967 \$9 dff_nclk
X$33469 \$1 \$9 \$I71961 \$I71962 \$I71964 \$I71963 sg13g2_or3_1
X$33470 \$I71962 \$41 \$I71960 \$I71966 \$I71969 \$1 \$I71961 \$9 freq_div_cell
X$33471 \$I71963 \$13 \$I71960 \$I71969 \$I71968 \$1 \$I71961 \$9 freq_div_cell
X$33472 \$9 \$1 \$I71968 sg13g2_tiehi
X$33473 \$I71964 \$48 \$I71960 \$I71970 \$I71966 \$1 \$I71961 \$9 freq_div_cell
M$1 \$1 \$42 \$I33319 \$1 sg13_lv_nmos L=0.13u W=1.2u AS=0.408p AD=0.228p
+ PS=3.08u PD=1.58u
M$2 \$I33319 \$10 \$43 \$1 sg13_lv_nmos L=0.13u W=1.2u AS=0.228p AD=0.408p
+ PS=1.58u PD=3.08u
M$3 \$43 \$I33318 \$46 \$9 sg13_lv_pmos L=0.13u W=0.15u AS=0.1005p AD=0.0555p
+ PS=1.34u PD=0.74u
M$4 \$46 \$45 \$9 \$9 sg13_lv_pmos L=0.13u W=0.15u AS=0.0555p AD=0.1005p
+ PS=0.74u PD=1.34u
M$5 \$25 \$23 \$22 \$1 sg13_lv_nmos L=0.13u W=1u AS=0.28p AD=0.28p PS=2.62u
+ PD=2.62u
M$7 \$1 \$28 \$I71937 \$1 sg13_lv_nmos L=0.13u W=0.6u AS=0.159p AD=0.159p
+ PS=1.96u PD=1.96u
M$9 \$1 \$28 \$26 \$1 sg13_lv_nmos L=0.13u W=0.6u AS=0.159p AD=0.159p PS=1.96u
+ PD=1.96u
M$11 \$1 \$28 \$I71939 \$1 sg13_lv_nmos L=0.13u W=0.6u AS=0.159p AD=0.159p
+ PS=1.96u PD=1.96u
M$13 \$1 \$28 \$I71940 \$1 sg13_lv_nmos L=0.13u W=0.6u AS=0.159p AD=0.159p
+ PS=1.96u PD=1.96u
M$15 \$26 \$21 \$20 \$1 sg13_lv_nmos L=0.13u W=1u AS=0.28p AD=0.28p PS=2.62u
+ PD=2.62u
M$17 \$1 \$28 \$I71941 \$1 sg13_lv_nmos L=0.13u W=0.6u AS=0.159p AD=0.159p
+ PS=1.96u PD=1.96u
M$19 \$I71936 \$24 \$23 \$1 sg13_lv_nmos L=0.13u W=1u AS=0.28p AD=0.28p
+ PS=2.62u PD=2.62u
M$21 \$I71935 \$22 \$21 \$1 sg13_lv_nmos L=0.13u W=1u AS=0.28p AD=0.28p
+ PS=2.62u PD=2.62u
M$23 \$I71937 \$8 \$24 \$1 sg13_lv_nmos L=0.13u W=1u AS=0.265p AD=0.265p
+ PS=2.56u PD=2.56u
M$25 \$1 \$28 \$I71935 \$1 sg13_lv_nmos L=0.13u W=0.6u AS=0.159p AD=0.159p
+ PS=1.96u PD=1.96u
M$27 \$1 \$28 \$25 \$1 sg13_lv_nmos L=0.13u W=0.6u AS=0.159p AD=0.159p PS=1.96u
+ PD=1.96u
M$29 \$1 \$28 \$I71942 \$1 sg13_lv_nmos L=0.13u W=0.6u AS=0.159p AD=0.159p
+ PS=1.96u PD=1.96u
M$31 \$1 \$28 \$I71938 \$1 sg13_lv_nmos L=0.13u W=0.6u AS=0.159p AD=0.159p
+ PS=1.96u PD=1.96u
M$33 \$1 \$28 \$14 \$1 sg13_lv_nmos L=0.13u W=0.6u AS=0.159p AD=0.159p PS=1.96u
+ PD=1.96u
M$35 \$1 \$28 \$I71934 \$1 sg13_lv_nmos L=0.13u W=0.6u AS=0.159p AD=0.159p
+ PS=1.96u PD=1.96u
M$37 \$1 \$28 \$I71936 \$1 sg13_lv_nmos L=0.13u W=0.6u AS=0.159p AD=0.159p
+ PS=1.96u PD=1.96u
M$39 \$I71934 \$20 \$I71933 \$1 sg13_lv_nmos L=0.13u W=1u AS=0.28p AD=0.28p
+ PS=2.62u PD=2.62u
M$41 \$9 \$14 \$I71927 \$9 sg13_lv_pmos L=0.13u W=0.8u AS=0.28325p AD=0.28175p
+ PS=3.575u PD=3.565u
M$45 \$I71930 \$8 \$24 \$9 sg13_lv_pmos L=0.13u W=2u AS=0.455p AD=0.455p
+ PS=4.32u PD=4.32u
M$49 \$9 \$14 \$14 \$9 sg13_lv_pmos L=0.13u W=0.8u AS=0.2825p AD=0.2825p
+ PS=3.57u PD=3.57u
M$53 \$9 \$14 \$I71945 \$9 sg13_lv_pmos L=0.13u W=0.8u AS=0.23825p AD=0.32675p
+ PS=2.975u PD=4.165u
M$57 \$9 \$14 \$I71931 \$9 sg13_lv_pmos L=0.13u W=0.8u AS=0.28325p AD=0.28175p
+ PS=3.575u PD=3.565u
M$61 \$9 \$14 \$I71944 \$9 sg13_lv_pmos L=0.13u W=0.8u AS=0.23825p AD=0.32675p
+ PS=2.975u PD=4.165u
M$65 \$I71929 \$24 \$23 \$9 sg13_lv_pmos L=0.13u W=2u AS=0.455p AD=0.455p
+ PS=4.32u PD=4.32u
M$69 \$I71931 \$20 \$I71933 \$9 sg13_lv_pmos L=0.13u W=2u AS=0.455p AD=0.455p
+ PS=4.32u PD=4.32u
M$73 \$9 \$14 \$I71928 \$9 sg13_lv_pmos L=0.13u W=0.8u AS=0.28325p AD=0.28175p
+ PS=3.575u PD=3.565u
M$77 \$I71927 \$22 \$21 \$9 sg13_lv_pmos L=0.13u W=2u AS=0.455p AD=0.455p
+ PS=4.32u PD=4.32u
M$81 \$I71932 \$21 \$20 \$9 sg13_lv_pmos L=0.13u W=2u AS=0.455p AD=0.455p
+ PS=4.32u PD=4.32u
M$85 \$9 \$14 \$I71929 \$9 sg13_lv_pmos L=0.13u W=0.8u AS=0.28325p AD=0.28175p
+ PS=3.575u PD=3.565u
M$89 \$9 \$14 \$I71930 \$9 sg13_lv_pmos L=0.13u W=0.8u AS=0.281p AD=0.281p
+ PS=3.56u PD=3.56u
M$93 \$9 \$14 \$I71932 \$9 sg13_lv_pmos L=0.13u W=0.8u AS=0.28325p AD=0.28175p
+ PS=3.575u PD=3.565u
M$97 \$9 \$14 \$I71946 \$9 sg13_lv_pmos L=0.13u W=0.8u AS=0.23825p AD=0.32675p
+ PS=2.975u PD=4.165u
M$101 \$9 \$14 \$I71943 \$9 sg13_lv_pmos L=0.13u W=0.8u AS=0.23825p AD=0.32675p
+ PS=2.975u PD=4.165u
M$105 \$9 \$14 \$I71947 \$9 sg13_lv_pmos L=0.13u W=0.8u AS=0.23825p AD=0.32675p
+ PS=2.975u PD=4.165u
M$109 \$I71928 \$23 \$22 \$9 sg13_lv_pmos L=0.13u W=2u AS=0.455p AD=0.455p
+ PS=4.32u PD=4.32u
M$113 \$I33318 \$44 \$9 \$9 sg13_lv_pmos L=0.13u W=0.3u AS=0.102p AD=0.102p
+ PS=1.28u PD=1.28u
M$114 \$1 \$44 \$I33318 \$1 sg13_lv_nmos L=0.13u W=0.15u AS=0.1005p AD=0.1005p
+ PS=1.34u PD=1.34u
C$115 \$21 \$1 cap_cmim w=6.99u l=6.99u A=48.8601p P=27.96u m=1
C$116 \$22 \$1 cap_cmim w=6.99u l=6.99u A=48.8601p P=27.96u m=1
C$117 \$31 \$1 cap_cmim w=6.99u l=6.99u A=48.8601p P=27.96u m=1
C$118 \$32 \$1 cap_cmim w=6.99u l=6.99u A=48.8601p P=27.96u m=1
C$119 \$I71933 \$1 cap_cmim w=6.99u l=6.99u A=48.8601p P=27.96u m=1
C$120 \$20 \$1 cap_cmim w=6.99u l=6.99u A=48.8601p P=27.96u m=1
C$121 \$23 \$1 cap_cmim w=6.99u l=6.99u A=48.8601p P=27.96u m=1
C$122 \$24 \$1 cap_cmim w=6.99u l=6.99u A=48.8601p P=27.96u m=1
C$123 \$34 \$1 cap_cmim w=6.99u l=6.99u A=48.8601p P=27.96u m=1
C$124 \$8 \$1 cap_cmim w=6.99u l=6.99u A=48.8601p P=27.96u m=1
C$125 \$33 \$1 cap_cmim w=6.99u l=6.99u A=48.8601p P=27.96u m=1
M$126 \$I71938 \$I71933 \$31 \$1 sg13_lv_nmos L=0.13u W=1u AS=0.265p AD=0.265p
+ PS=2.56u PD=2.56u
M$128 \$I71943 \$I71933 \$31 \$9 sg13_lv_pmos L=0.13u W=2u AS=0.455p AD=0.455p
+ PS=4.32u PD=4.32u
M$132 \$I71939 \$31 \$32 \$1 sg13_lv_nmos L=0.13u W=1u AS=0.265p AD=0.265p
+ PS=2.56u PD=2.56u
M$134 \$I71944 \$31 \$32 \$9 sg13_lv_pmos L=0.13u W=2u AS=0.455p AD=0.455p
+ PS=4.32u PD=4.32u
M$138 \$I71941 \$32 \$33 \$1 sg13_lv_nmos L=0.13u W=1u AS=0.265p AD=0.265p
+ PS=2.56u PD=2.56u
M$140 \$I71945 \$32 \$33 \$9 sg13_lv_pmos L=0.13u W=2u AS=0.455p AD=0.455p
+ PS=4.32u PD=4.32u
M$144 \$I71942 \$33 \$34 \$1 sg13_lv_nmos L=0.13u W=1u AS=0.265p AD=0.265p
+ PS=2.56u PD=2.56u
M$146 \$I71946 \$33 \$34 \$9 sg13_lv_pmos L=0.13u W=2u AS=0.455p AD=0.455p
+ PS=4.32u PD=4.32u
M$150 \$I71940 \$34 \$8 \$1 sg13_lv_nmos L=0.13u W=1u AS=0.265p AD=0.265p
+ PS=2.56u PD=2.56u
M$152 \$I71947 \$34 \$8 \$9 sg13_lv_pmos L=0.13u W=2u AS=0.455p AD=0.455p
+ PS=4.32u PD=4.32u
.ENDS FMD_QNC_PLL_3BIT_DIV

.SUBCKT PFD VDD VSS DOWN VCO_CLK UP Ref_CLK
M$1 \$5 VCO_CLK \$7 VSS sg13_lv_nmos L=0.15u W=0.84u AS=0.2226p AD=0.2226p
+ PS=2.32u PD=2.32u
M$3 \$10 Ref_CLK \$12 VSS sg13_lv_nmos L=0.15u W=0.84u AS=0.2226p AD=0.2226p
+ PS=2.32u PD=2.32u
M$5 VSS \$13 UP VSS sg13_lv_nmos L=0.15u W=0.48u AS=0.1632p AD=0.1632p PS=1.64u
+ PD=1.64u
M$6 VSS \$4 DOWN VSS sg13_lv_nmos L=0.15u W=0.48u AS=0.1632p AD=0.1632p
+ PS=1.64u PD=1.64u
M$7 \$8 VCO_CLK VSS VSS sg13_lv_nmos L=0.15u W=0.36u AS=0.1224p AD=0.1224p
+ PS=1.4u PD=1.4u
M$8 VSS \$10 \$13 VSS sg13_lv_nmos L=0.15u W=0.36u AS=0.1224p AD=0.1224p
+ PS=1.4u PD=1.4u
M$9 VSS \$5 \$4 VSS sg13_lv_nmos L=0.15u W=0.36u AS=0.1224p AD=0.1224p PS=1.4u
+ PD=1.4u
M$10 \$9 Ref_CLK VSS VSS sg13_lv_nmos L=0.15u W=0.36u AS=0.1224p AD=0.1224p
+ PS=1.4u PD=1.4u
M$11 VDD \$13 UP VDD sg13_lv_pmos L=0.15u W=0.96u AS=0.2304p AD=0.2304p
+ PS=2.72u PD=2.72u
M$14 VDD \$4 DOWN VDD sg13_lv_pmos L=0.15u W=0.96u AS=0.2304p AD=0.2304p
+ PS=2.72u PD=2.72u
M$17 \$13 \$10 VDD VDD sg13_lv_pmos L=0.15u W=0.72u AS=0.1908p AD=0.1908p
+ PS=2.14u PD=2.14u
M$19 VDD \$5 \$4 VDD sg13_lv_pmos L=0.15u W=0.72u AS=0.1908p AD=0.1908p
+ PS=2.14u PD=2.14u
M$21 \$8 Ref_CLK \$12 VSS sg13_lv_nmos L=0.15u W=1.8u AS=0.396p AD=0.396p
+ PS=4.36u PD=4.36u
M$26 \$9 VCO_CLK \$7 VSS sg13_lv_nmos L=0.15u W=1.8u AS=0.396p AD=0.396p
+ PS=4.36u PD=4.36u
M$31 \$12 Ref_CLK VDD VDD sg13_lv_pmos L=0.15u W=0.64u AS=0.1696p AD=0.1696p
+ PS=2.02u PD=2.02u
M$33 \$7 VCO_CLK VDD VDD sg13_lv_pmos L=0.15u W=0.64u AS=0.1696p AD=0.1696p
+ PS=2.02u PD=2.02u
M$35 \$5 VCO_CLK VCO_CLK VDD sg13_lv_pmos L=0.15u W=0.64u AS=0.1696p AD=0.1696p
+ PS=2.02u PD=2.02u
M$37 \$10 Ref_CLK Ref_CLK VDD sg13_lv_pmos L=0.15u W=0.64u AS=0.1696p
+ AD=0.1696p PS=2.02u PD=2.02u
.ENDS PFD

.SUBCKT Bias_gen \$1 \$2 enb en \$6 \$9 \$10 \$13
R$1 \$11 \$13 rhigh w=1u l=12u ps=0 b=0 m=1
R$2 \$3 \$2 rhigh w=1u l=12u ps=0 b=0 m=1
M$3 \$7 \$6 \$2 \$1 sg13_lv_nmos L=1u W=1u AS=0.34p AD=0.34p PS=2.68u PD=2.68u
M$4 \$9 \$6 \$3 \$1 sg13_lv_nmos L=1u W=1u AS=0.34p AD=0.34p PS=2.68u PD=2.68u
M$5 \$6 \$6 \$2 \$1 sg13_lv_nmos L=1u W=1u AS=0.34p AD=0.34p PS=2.68u PD=2.68u
M$6 \$9 \$7 \$8 \$1 sg13_lv_nmos L=0.15u W=0.5u AS=0.17p AD=0.17p PS=1.68u
+ PD=1.68u
M$7 \$6 enb \$2 \$1 sg13_lv_nmos L=0.15u W=0.5u AS=0.17p AD=0.17p PS=1.68u
+ PD=1.68u
M$8 \$8 en \$2 \$1 sg13_lv_nmos L=0.15u W=0.5u AS=0.17p AD=0.17p PS=1.68u
+ PD=1.68u
M$9 \$6 \$9 \$11 \$10 sg13_lv_pmos L=1u W=4u AS=1.06p AD=1.06p PS=7.06u PD=7.06u
M$11 \$13 \$9 \$9 \$10 sg13_lv_pmos L=1u W=2u AS=0.68p AD=0.68p PS=4.68u
+ PD=4.68u
M$12 \$13 \$12 \$12 \$10 sg13_lv_pmos L=0.15u W=0.5u AS=0.17p AD=0.17p PS=1.68u
+ PD=1.68u
M$13 \$13 en \$9 \$10 sg13_lv_pmos L=0.15u W=0.5u AS=0.17p AD=0.17p PS=1.68u
+ PD=1.68u
M$14 \$12 \$7 \$7 \$10 sg13_lv_pmos L=0.15u W=0.5u AS=0.17p AD=0.17p PS=1.68u
+ PD=1.68u
M$15 \$13 en \$7 \$10 sg13_lv_pmos L=0.15u W=0.5u AS=0.17p AD=0.17p PS=1.68u
+ PD=1.68u
.ENDS Bias_gen

.SUBCKT loop_filter \$1 \$2 \$3
M$1 \$1 \$2 \$1 \$1 sg13_lv_nmos L=0.65u W=45u AS=9p AD=9p PS=60u PD=60u
R$31 \$2 \$3 rhigh w=0.6u l=0.96u ps=0 b=0 m=1
R$32 \$4 \$2 rhigh w=0.5u l=0.96u ps=0 b=0 m=1
M$33 \$1 \$3 \$1 \$1 sg13_lv_nmos L=0.13u W=0.3u AS=0.201p AD=0.201p PS=2.68u
+ PD=2.68u
M$35 \$1 \$4 \$1 \$1 sg13_lv_nmos L=0.65u W=15u AS=3p AD=3p PS=28u PD=28u
.ENDS loop_filter

.SUBCKT sg13g2_nand2_1 VSS VDD Y B A
M$1 VSS B \$6 VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.2516p AD=0.0666p PS=2.16u
+ PD=0.92u
M$2 \$6 A Y VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.0666p AD=0.2516p PS=0.92u
+ PD=2.16u
M$3 VDD B Y VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.3808p AD=0.2128p PS=2.92u
+ PD=1.5u
M$4 Y A VDD VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.2128p AD=0.3808p PS=1.5u
+ PD=2.92u
.ENDS sg13g2_nand2_1

.SUBCKT sg13g2_or3_1 VSS VDD X B A C
M$1 \$4 C VSS VSS sg13_lv_nmos L=0.13u W=0.55u AS=0.187p AD=0.1045p PS=1.78u
+ PD=0.93u
M$2 VSS B \$4 VSS sg13_lv_nmos L=0.13u W=0.55u AS=0.1045p AD=0.198p PS=0.93u
+ PD=1.27u
M$3 \$4 A VSS VSS sg13_lv_nmos L=0.13u W=0.55u AS=0.198p AD=0.13395p PS=1.27u
+ PD=1.12u
M$4 VSS \$4 X VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.13395p AD=0.2516p PS=1.12u
+ PD=2.16u
M$5 \$4 C \$9 VDD sg13_lv_pmos L=0.13u W=1u AS=0.34p AD=0.1275p PS=2.68u
+ PD=1.255u
M$6 \$9 B \$8 VDD sg13_lv_pmos L=0.13u W=1u AS=0.1275p AD=0.22p PS=1.255u
+ PD=1.44u
M$7 \$8 A VDD VDD sg13_lv_pmos L=0.13u W=1u AS=0.22p AD=0.3822p PS=1.44u
+ PD=1.84u
M$8 VDD \$4 X VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.3822p AD=0.3808p PS=1.84u
+ PD=2.92u
.ENDS sg13g2_or3_1

.SUBCKT sg13g2_tiehi VDD VSS L_HI
M$1 VSS \$3 \$3 VSS sg13_lv_nmos L=0.13u W=0.3u AS=0.2307p AD=0.102p PS=1.615u
+ PD=1.28u
M$2 VSS \$4 \$6 VSS sg13_lv_nmos L=0.13u W=0.795u AS=0.2307p AD=0.274275p
+ PS=1.615u PD=2.28u
M$3 \$4 \$3 VDD VDD sg13_lv_pmos L=0.13u W=0.66u AS=0.2442p AD=0.4657125p
+ PS=2.06u PD=2.54u
M$4 VDD \$6 L_HI VDD sg13_lv_pmos L=0.13u W=1.155u AS=0.4657125p AD=0.3927p
+ PS=2.54u PD=2.99u
.ENDS sg13g2_tiehi

.SUBCKT freq_div_cell DIV BIT CLK Cout Cin \$7 nRST \$12
X$1 BIT \$12 DIV \$7 \$6 sg13g2_xor2_1
X$2 \$6 \$I8 \$8 CLK \$7 nRST \$12 dff_nclk
X$3 Cout \$8 \$6 Cin \$7 \$12 half_add
.ENDS freq_div_cell

.SUBCKT dff_nclk Q nQ D nCLK \$6 nRST \$8
X$1 \$6 nRST nQ Q D \$5 \$8 sg13g2_dfrbp_1
X$2 \$8 \$6 nCLK \$5 sg13g2_inv_1
.ENDS dff_nclk

.SUBCKT half_add cout sum inB inA \$5 \$7
X$1 \$7 \$5 cout inB inA sg13g2_and2_1
X$2 inB \$7 sum \$5 inA sg13g2_xor2_1
.ENDS half_add

.SUBCKT sg13g2_dfrbp_1 VSS RESET_B Q_N Q D CLK VDD
M$1 \$5 \$11 \$19 VSS sg13_lv_nmos L=0.13u W=0.42u AS=0.2017p AD=0.0546p
+ PS=1.48u PD=0.68u
M$2 \$19 \$6 VSS VSS sg13_lv_nmos L=0.13u W=0.42u AS=0.0546p AD=0.0903p
+ PS=0.68u PD=0.85u
M$3 VSS RESET_B \$18 VSS sg13_lv_nmos L=0.13u W=0.42u AS=0.0903p AD=0.04725p
+ PS=0.85u PD=0.645u
M$4 \$18 \$5 \$6 VSS sg13_lv_nmos L=0.13u W=0.42u AS=0.04725p AD=0.1428p
+ PS=0.645u PD=1.52u
M$5 VSS \$13 \$14 VSS sg13_lv_nmos L=0.13u W=0.64u AS=0.1825p AD=0.193975p
+ PS=1.325u PD=1.29u
M$6 \$14 \$3 \$5 VSS sg13_lv_nmos L=0.13u W=0.64u AS=0.193975p AD=0.2017p
+ PS=1.29u PD=1.48u
M$7 \$4 \$11 \$13 VSS sg13_lv_nmos L=0.13u W=0.42u AS=0.1428p AD=0.0798p
+ PS=1.52u PD=0.8u
M$8 \$13 \$3 \$16 VSS sg13_lv_nmos L=0.13u W=0.42u AS=0.0798p AD=0.0546p
+ PS=0.8u PD=0.68u
M$9 \$16 \$14 \$17 VSS sg13_lv_nmos L=0.13u W=0.42u AS=0.0546p AD=0.0483p
+ PS=0.68u PD=0.65u
M$10 VSS RESET_B \$17 VSS sg13_lv_nmos L=0.13u W=0.42u AS=0.1825p AD=0.0483p
+ PS=1.325u PD=0.65u
M$11 \$8 \$5 VSS VSS sg13_lv_nmos L=0.13u W=0.55u AS=0.187p AD=0.14505p
+ PS=1.78u PD=1.15u
M$12 VSS \$8 Q VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.14505p AD=0.2516p PS=1.15u
+ PD=2.16u
M$13 VSS \$5 Q_N VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.2516p AD=0.2775p
+ PS=2.16u PD=2.23u
M$14 VSS CLK \$11 VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.1544p AD=0.2516p
+ PS=1.235u PD=2.16u
M$15 VSS \$11 \$3 VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.1544p AD=0.2516p
+ PS=1.235u PD=2.16u
M$16 \$4 D \$15 VSS sg13_lv_nmos L=0.13u W=0.42u AS=0.1428p AD=0.0504p PS=1.52u
+ PD=0.66u
M$17 \$15 RESET_B VSS VSS sg13_lv_nmos L=0.13u W=0.42u AS=0.0504p AD=0.1428p
+ PS=0.66u PD=1.52u
M$18 VDD \$13 \$14 VDD sg13_lv_pmos L=0.13u W=1u AS=0.34p AD=0.19p PS=2.68u
+ PD=1.38u
M$19 \$14 \$11 \$5 VDD sg13_lv_pmos L=0.13u W=1u AS=0.19p AD=0.17695p PS=1.38u
+ PD=1.56u
M$20 \$5 \$3 \$22 VDD sg13_lv_pmos L=0.13u W=0.42u AS=0.17695p AD=0.04305p
+ PS=1.56u PD=0.625u
M$21 \$22 \$6 VDD VDD sg13_lv_pmos L=0.13u W=0.42u AS=0.04305p AD=0.0798p
+ PS=0.625u PD=0.8u
M$22 VDD RESET_B \$6 VDD sg13_lv_pmos L=0.13u W=0.42u AS=0.0798p AD=0.0798p
+ PS=0.8u PD=0.8u
M$23 VDD \$5 \$6 VDD sg13_lv_pmos L=0.13u W=0.42u AS=0.2163p AD=0.0798p
+ PS=1.55u PD=0.8u
M$24 VDD \$5 Q_N VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.2163p AD=0.7616p
+ PS=1.55u PD=3.6u
M$25 \$4 \$3 \$13 VDD sg13_lv_pmos L=0.13u W=0.42u AS=0.1428p AD=0.0798p
+ PS=1.52u PD=0.8u
M$26 \$13 \$11 \$21 VDD sg13_lv_pmos L=0.13u W=0.42u AS=0.0798p AD=0.05145p
+ PS=0.8u PD=0.665u
M$27 \$21 \$14 VDD VDD sg13_lv_pmos L=0.13u W=0.42u AS=0.05145p AD=0.11785p
+ PS=0.665u PD=1.025u
M$28 VDD RESET_B \$13 VDD sg13_lv_pmos L=0.13u W=0.42u AS=0.11785p AD=0.1533p
+ PS=1.025u PD=1.57u
M$29 \$11 CLK VDD VDD sg13_lv_pmos L=0.13u W=1u AS=0.34p AD=0.19p PS=2.68u
+ PD=1.38u
M$30 VDD \$11 \$3 VDD sg13_lv_pmos L=0.13u W=1u AS=0.19p AD=0.34p PS=1.38u
+ PD=2.68u
M$31 VDD D \$4 VDD sg13_lv_pmos L=0.13u W=0.42u AS=0.1428p AD=0.0798p PS=1.52u
+ PD=0.8u
M$32 \$4 RESET_B VDD VDD sg13_lv_pmos L=0.13u W=0.42u AS=0.0798p AD=0.1428p
+ PS=0.8u PD=1.52u
M$33 VDD \$5 \$8 VDD sg13_lv_pmos L=0.13u W=0.84u AS=0.2016p AD=0.2856p PS=1.5u
+ PD=2.36u
M$34 VDD \$8 Q VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.2016p AD=0.3808p PS=1.5u
+ PD=2.92u
.ENDS sg13g2_dfrbp_1

.SUBCKT sg13g2_inv_1 VDD VSS A Y
M$1 VSS A Y VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.259p AD=0.259p PS=2.18u
+ PD=2.18u
M$2 VDD A Y VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.392p AD=0.392p PS=2.94u
+ PD=2.94u
.ENDS sg13g2_inv_1

.SUBCKT sg13g2_and2_1 VDD VSS X B A
M$1 \$3 A \$7 VSS sg13_lv_nmos L=0.13u W=0.64u AS=0.2176p AD=0.1216p PS=1.96u
+ PD=1.02u
M$2 VSS B \$7 VSS sg13_lv_nmos L=0.13u W=0.64u AS=0.1331p AD=0.1216p PS=1.12u
+ PD=1.02u
M$3 VSS \$3 X VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.1331p AD=0.2516p PS=1.12u
+ PD=2.16u
M$4 VDD A \$3 VDD sg13_lv_pmos L=0.13u W=0.84u AS=0.2856p AD=0.1596p PS=2.36u
+ PD=1.22u
M$5 VDD B \$3 VDD sg13_lv_pmos L=0.13u W=0.84u AS=0.1918p AD=0.1596p PS=1.5u
+ PD=1.22u
M$6 VDD \$3 X VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.1918p AD=0.3808p PS=1.5u
+ PD=2.92u
.ENDS sg13g2_and2_1

.SUBCKT sg13g2_xor2_1 B VDD X VSS A
M$1 VSS A \$7 VSS sg13_lv_nmos L=0.13u W=0.55u AS=0.374p AD=0.174625p PS=2.46u
+ PD=1.185u
M$2 VSS B \$7 VSS sg13_lv_nmos L=0.13u W=0.55u AS=0.15245p AD=0.174625p
+ PS=1.17u PD=1.185u
M$3 VSS A \$8 VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.15245p AD=0.0888p PS=1.17u
+ PD=0.98u
M$4 \$8 B X VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.0888p AD=0.1628p PS=0.98u
+ PD=1.18u
M$5 X \$7 VSS VSS sg13_lv_nmos L=0.13u W=0.74u AS=0.1628p AD=0.3108p PS=1.18u
+ PD=2.32u
M$6 \$2 A VDD VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.3808p AD=0.2128p PS=2.92u
+ PD=1.5u
M$7 VDD B \$2 VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.2128p AD=0.2128p PS=1.5u
+ PD=1.5u
M$8 \$2 \$7 X VDD sg13_lv_pmos L=0.13u W=1.12u AS=0.2128p AD=0.3808p PS=1.5u
+ PD=2.92u
M$9 VDD A \$9 VDD sg13_lv_pmos L=0.13u W=1u AS=0.36p AD=0.1225p PS=2.72u
+ PD=1.245u
M$10 \$9 B \$7 VDD sg13_lv_pmos L=0.13u W=1u AS=0.1225p AD=0.34p PS=1.245u
+ PD=2.68u
.ENDS sg13g2_xor2_1
